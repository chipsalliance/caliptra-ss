// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef MCI_REG_DEFINES_HEADER
`define MCI_REG_DEFINES_HEADER


`define MCI_REG_BASE_ADDR                                                                           (32'h0)
`define MCI_REG_CAPABILITIES                                                                        (32'h0)
`define MCI_REG_CAPABILITIES                                                                        (32'h0)
`define MCI_REG_CAPABILITIES_NUM_MBOX_LOW                                                           (0)
`define MCI_REG_CAPABILITIES_NUM_MBOX_MASK                                                          (32'hf)
`define MCI_REG_HW_REV_ID                                                                           (32'h4)
`define MCI_REG_HW_REV_ID                                                                           (32'h4)
`define MCI_REG_HW_REV_ID_MC_GENERATION_LOW                                                         (0)
`define MCI_REG_HW_REV_ID_MC_GENERATION_MASK                                                        (32'hffff)
`define MCI_REG_HW_REV_ID_SOC_STEPPING_ID_LOW                                                       (16)
`define MCI_REG_HW_REV_ID_SOC_STEPPING_ID_MASK                                                      (32'hffff0000)
`define MCI_REG_FW_REV_ID_0                                                                         (32'h8)
`define MCI_REG_FW_REV_ID_0                                                                         (32'h8)
`define MCI_REG_FW_REV_ID_1                                                                         (32'hc)
`define MCI_REG_FW_REV_ID_1                                                                         (32'hc)
`define MCI_REG_HW_CONFIG                                                                           (32'h10)
`define MCI_REG_HW_CONFIG                                                                           (32'h10)
`define MCI_REG_HW_CONFIG_RSVD_EN_LOW                                                               (0)
`define MCI_REG_HW_CONFIG_RSVD_EN_MASK                                                              (32'h1)
`define MCI_REG_FW_FLOW_STATUS                                                                      (32'h20)
`define MCI_REG_FW_FLOW_STATUS                                                                      (32'h20)
`define MCI_REG_HW_FLOW_STATUS                                                                      (32'h24)
`define MCI_REG_HW_FLOW_STATUS                                                                      (32'h24)
`define MCI_REG_HW_FLOW_STATUS_BOOT_FSM_LOW                                                         (0)
`define MCI_REG_HW_FLOW_STATUS_BOOT_FSM_MASK                                                        (32'hf)
`define MCI_REG_RESET_REASON                                                                        (32'h28)
`define MCI_REG_RESET_REASON                                                                        (32'h28)
`define MCI_REG_RESET_REASON_FW_HITLESS_UPD_RESET_LOW                                               (0)
`define MCI_REG_RESET_REASON_FW_HITLESS_UPD_RESET_MASK                                              (32'h1)
`define MCI_REG_RESET_REASON_FW_BOOT_UPD_RESET_LOW                                                  (1)
`define MCI_REG_RESET_REASON_FW_BOOT_UPD_RESET_MASK                                                 (32'h2)
`define MCI_REG_RESET_REASON_WARM_RESET_LOW                                                         (2)
`define MCI_REG_RESET_REASON_WARM_RESET_MASK                                                        (32'h4)
`define MCI_REG_RESET_STATUS                                                                        (32'h2c)
`define MCI_REG_RESET_STATUS                                                                        (32'h2c)
`define MCI_REG_RESET_STATUS_CPTRA_RESET_STS_LOW                                                    (0)
`define MCI_REG_RESET_STATUS_CPTRA_RESET_STS_MASK                                                   (32'h1)
`define MCI_REG_RESET_STATUS_MCU_RESET_STS_LOW                                                      (1)
`define MCI_REG_RESET_STATUS_MCU_RESET_STS_MASK                                                     (32'h2)
`define MCI_REG_HW_ERROR_FATAL                                                                      (32'h40)
`define MCI_REG_HW_ERROR_FATAL                                                                      (32'h40)
`define MCI_REG_HW_ERROR_FATAL_MCU_SRAM_ECC_UNC_LOW                                                 (0)
`define MCI_REG_HW_ERROR_FATAL_MCU_SRAM_ECC_UNC_MASK                                                (32'h1)
`define MCI_REG_HW_ERROR_FATAL_NMI_PIN_LOW                                                          (1)
`define MCI_REG_HW_ERROR_FATAL_NMI_PIN_MASK                                                         (32'h2)
`define MCI_REG_AGG_ERROR_FATAL                                                                     (32'h44)
`define MCI_REG_AGG_ERROR_FATAL                                                                     (32'h44)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL31_LOW                                               (0)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL31_MASK                                              (32'h1)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL30_LOW                                               (1)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL30_MASK                                              (32'h2)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL29_LOW                                               (2)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL29_MASK                                              (32'h4)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL28_LOW                                               (3)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL28_MASK                                              (32'h8)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL27_LOW                                               (4)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL27_MASK                                              (32'h10)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL26_LOW                                               (5)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL26_MASK                                              (32'h20)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL25_LOW                                               (6)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL25_MASK                                              (32'h40)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL24_LOW                                               (7)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL24_MASK                                              (32'h80)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL23_LOW                                               (8)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL23_MASK                                              (32'h100)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL22_LOW                                               (9)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL22_MASK                                              (32'h200)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL21_LOW                                               (10)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL21_MASK                                              (32'h400)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL20_LOW                                               (11)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL20_MASK                                              (32'h800)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL19_LOW                                               (12)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL19_MASK                                              (32'h1000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL18_LOW                                               (13)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL18_MASK                                              (32'h2000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL17_LOW                                               (14)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL17_MASK                                              (32'h4000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL16_LOW                                               (15)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL16_MASK                                              (32'h8000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL15_LOW                                               (16)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL15_MASK                                              (32'h10000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL14_LOW                                               (17)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL14_MASK                                              (32'h20000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL13_LOW                                               (18)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL13_MASK                                              (32'h40000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL12_LOW                                               (19)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL12_MASK                                              (32'h80000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL11_LOW                                               (20)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL11_MASK                                              (32'h100000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL10_LOW                                               (21)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL10_MASK                                              (32'h200000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL9_LOW                                                (22)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL9_MASK                                               (32'h400000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL8_LOW                                                (23)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL8_MASK                                               (32'h800000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL7_LOW                                                (24)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL7_MASK                                               (32'h1000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL6_LOW                                                (25)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL6_MASK                                               (32'h2000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL5_LOW                                                (26)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL5_MASK                                               (32'h4000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL4_LOW                                                (27)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL4_MASK                                               (32'h8000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL3_LOW                                                (28)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL3_MASK                                               (32'h10000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL2_LOW                                                (29)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL2_MASK                                               (32'h20000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL1_LOW                                                (30)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL1_MASK                                               (32'h40000000)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL0_LOW                                                (31)
`define MCI_REG_AGG_ERROR_FATAL_AGG_ERROR_FATAL0_MASK                                               (32'h80000000)
`define MCI_REG_HW_ERROR_NON_FATAL                                                                  (32'h48)
`define MCI_REG_HW_ERROR_NON_FATAL                                                                  (32'h48)
`define MCI_REG_HW_ERROR_NON_FATAL_RSVD_LOW                                                         (0)
`define MCI_REG_HW_ERROR_NON_FATAL_RSVD_MASK                                                        (32'h1)
`define MCI_REG_AGG_ERROR_NON_FATAL                                                                 (32'h4c)
`define MCI_REG_AGG_ERROR_NON_FATAL                                                                 (32'h4c)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL31_LOW                                       (0)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL31_MASK                                      (32'h1)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL30_LOW                                       (1)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL30_MASK                                      (32'h2)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL29_LOW                                       (2)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL29_MASK                                      (32'h4)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL28_LOW                                       (3)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL28_MASK                                      (32'h8)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL27_LOW                                       (4)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL27_MASK                                      (32'h10)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL26_LOW                                       (5)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL26_MASK                                      (32'h20)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL25_LOW                                       (6)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL25_MASK                                      (32'h40)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL24_LOW                                       (7)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL24_MASK                                      (32'h80)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL23_LOW                                       (8)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL23_MASK                                      (32'h100)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL22_LOW                                       (9)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL22_MASK                                      (32'h200)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL21_LOW                                       (10)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL21_MASK                                      (32'h400)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL20_LOW                                       (11)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL20_MASK                                      (32'h800)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL19_LOW                                       (12)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL19_MASK                                      (32'h1000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL18_LOW                                       (13)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL18_MASK                                      (32'h2000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL17_LOW                                       (14)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL17_MASK                                      (32'h4000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL16_LOW                                       (15)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL16_MASK                                      (32'h8000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL15_LOW                                       (16)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL15_MASK                                      (32'h10000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL14_LOW                                       (17)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL14_MASK                                      (32'h20000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL13_LOW                                       (18)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL13_MASK                                      (32'h40000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL12_LOW                                       (19)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL12_MASK                                      (32'h80000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL11_LOW                                       (20)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL11_MASK                                      (32'h100000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL10_LOW                                       (21)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL10_MASK                                      (32'h200000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL9_LOW                                        (22)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL9_MASK                                       (32'h400000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL8_LOW                                        (23)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL8_MASK                                       (32'h800000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL7_LOW                                        (24)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL7_MASK                                       (32'h1000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL6_LOW                                        (25)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL6_MASK                                       (32'h2000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL5_LOW                                        (26)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL5_MASK                                       (32'h4000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL4_LOW                                        (27)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL4_MASK                                       (32'h8000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL3_LOW                                        (28)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL3_MASK                                       (32'h10000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL2_LOW                                        (29)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL2_MASK                                       (32'h20000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL1_LOW                                        (30)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL1_MASK                                       (32'h40000000)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL0_LOW                                        (31)
`define MCI_REG_AGG_ERROR_NON_FATAL_AGG_ERROR_NON_FATAL0_MASK                                       (32'h80000000)
`define MCI_REG_FW_ERROR_FATAL                                                                      (32'h50)
`define MCI_REG_FW_ERROR_FATAL                                                                      (32'h50)
`define MCI_REG_FW_ERROR_NON_FATAL                                                                  (32'h54)
`define MCI_REG_FW_ERROR_NON_FATAL                                                                  (32'h54)
`define MCI_REG_HW_ERROR_ENC                                                                        (32'h58)
`define MCI_REG_HW_ERROR_ENC                                                                        (32'h58)
`define MCI_REG_FW_ERROR_ENC                                                                        (32'h5c)
`define MCI_REG_FW_ERROR_ENC                                                                        (32'h5c)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_0                                                            (32'h60)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_0                                                            (32'h60)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_1                                                            (32'h64)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_1                                                            (32'h64)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_2                                                            (32'h68)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_2                                                            (32'h68)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_3                                                            (32'h6c)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_3                                                            (32'h6c)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_4                                                            (32'h70)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_4                                                            (32'h70)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_5                                                            (32'h74)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_5                                                            (32'h74)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_6                                                            (32'h78)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_6                                                            (32'h78)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_7                                                            (32'h7c)
`define MCI_REG_FW_EXTENDED_ERROR_INFO_7                                                            (32'h7c)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                        (32'h80)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                        (32'h80)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_MCU_SRAM_ECC_UNC_LOW                              (0)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_MCU_SRAM_ECC_UNC_MASK                             (32'h1)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_NMI_PIN_LOW                                       (1)
`define MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_NMI_PIN_MASK                                      (32'h2)
`define MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                                    (32'h84)
`define MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                                    (32'h84)
`define MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_FIXME_LOW                                          (0)
`define MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_FIXME_MASK                                         (32'h1)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK                                                       (32'h88)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK                                                       (32'h88)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL31_LOW                            (0)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL31_MASK                           (32'h1)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL30_LOW                            (1)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL30_MASK                           (32'h2)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL29_LOW                            (2)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL29_MASK                           (32'h4)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL28_LOW                            (3)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL28_MASK                           (32'h8)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL27_LOW                            (4)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL27_MASK                           (32'h10)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL26_LOW                            (5)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL26_MASK                           (32'h20)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL25_LOW                            (6)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL25_MASK                           (32'h40)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL24_LOW                            (7)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL24_MASK                           (32'h80)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL23_LOW                            (8)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL23_MASK                           (32'h100)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL22_LOW                            (9)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL22_MASK                           (32'h200)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL21_LOW                            (10)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL21_MASK                           (32'h400)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL20_LOW                            (11)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL20_MASK                           (32'h800)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL19_LOW                            (12)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL19_MASK                           (32'h1000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL18_LOW                            (13)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL18_MASK                           (32'h2000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL17_LOW                            (14)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL17_MASK                           (32'h4000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL16_LOW                            (15)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL16_MASK                           (32'h8000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL15_LOW                            (16)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL15_MASK                           (32'h10000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL14_LOW                            (17)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL14_MASK                           (32'h20000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL13_LOW                            (18)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL13_MASK                           (32'h40000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL12_LOW                            (19)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL12_MASK                           (32'h80000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL11_LOW                            (20)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL11_MASK                           (32'h100000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL10_LOW                            (21)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL10_MASK                           (32'h200000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL9_LOW                             (22)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL9_MASK                            (32'h400000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL8_LOW                             (23)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL8_MASK                            (32'h800000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL7_LOW                             (24)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL7_MASK                            (32'h1000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL6_LOW                             (25)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL6_MASK                            (32'h2000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL5_LOW                             (26)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL5_MASK                            (32'h4000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL4_LOW                             (27)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL4_MASK                            (32'h8000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL3_LOW                             (28)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL3_MASK                            (32'h10000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL2_LOW                             (29)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL2_MASK                            (32'h20000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL1_LOW                             (30)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL1_MASK                            (32'h40000000)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL0_LOW                             (31)
`define MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK_MASK_AGG_ERROR_FATAL0_MASK                            (32'h80000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK                                                   (32'h8c)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK                                                   (32'h8c)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL31_LOW                    (0)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL31_MASK                   (32'h1)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL30_LOW                    (1)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL30_MASK                   (32'h2)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL29_LOW                    (2)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL29_MASK                   (32'h4)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL28_LOW                    (3)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL28_MASK                   (32'h8)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL27_LOW                    (4)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL27_MASK                   (32'h10)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL26_LOW                    (5)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL26_MASK                   (32'h20)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL25_LOW                    (6)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL25_MASK                   (32'h40)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL24_LOW                    (7)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL24_MASK                   (32'h80)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL23_LOW                    (8)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL23_MASK                   (32'h100)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL22_LOW                    (9)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL22_MASK                   (32'h200)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL21_LOW                    (10)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL21_MASK                   (32'h400)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL20_LOW                    (11)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL20_MASK                   (32'h800)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL19_LOW                    (12)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL19_MASK                   (32'h1000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL18_LOW                    (13)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL18_MASK                   (32'h2000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL17_LOW                    (14)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL17_MASK                   (32'h4000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL16_LOW                    (15)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL16_MASK                   (32'h8000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL15_LOW                    (16)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL15_MASK                   (32'h10000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL14_LOW                    (17)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL14_MASK                   (32'h20000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL13_LOW                    (18)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL13_MASK                   (32'h40000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL12_LOW                    (19)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL12_MASK                   (32'h80000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL11_LOW                    (20)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL11_MASK                   (32'h100000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL10_LOW                    (21)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL10_MASK                   (32'h200000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL9_LOW                     (22)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL9_MASK                    (32'h400000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL8_LOW                     (23)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL8_MASK                    (32'h800000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL7_LOW                     (24)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL7_MASK                    (32'h1000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL6_LOW                     (25)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL6_MASK                    (32'h2000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL5_LOW                     (26)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL5_MASK                    (32'h4000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL4_LOW                     (27)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL4_MASK                    (32'h8000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL3_LOW                     (28)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL3_MASK                    (32'h10000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL2_LOW                     (29)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL2_MASK                    (32'h20000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL1_LOW                     (30)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL1_MASK                    (32'h40000000)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL0_LOW                     (31)
`define MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK_MASK_AGG_ERROR_NON_FATAL0_MASK                    (32'h80000000)
`define MCI_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                        (32'h90)
`define MCI_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                        (32'h90)
`define MCI_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                                    (32'h94)
`define MCI_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                                    (32'h94)
`define MCI_REG_WDT_TIMER1_EN                                                                       (32'ha0)
`define MCI_REG_WDT_TIMER1_EN                                                                       (32'ha0)
`define MCI_REG_WDT_TIMER1_EN_TIMER1_EN_LOW                                                         (0)
`define MCI_REG_WDT_TIMER1_EN_TIMER1_EN_MASK                                                        (32'h1)
`define MCI_REG_WDT_TIMER1_CTRL                                                                     (32'ha4)
`define MCI_REG_WDT_TIMER1_CTRL                                                                     (32'ha4)
`define MCI_REG_WDT_TIMER1_CTRL_TIMER1_RESTART_LOW                                                  (0)
`define MCI_REG_WDT_TIMER1_CTRL_TIMER1_RESTART_MASK                                                 (32'h1)
`define MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_0                                                         (32'ha8)
`define MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_0                                                         (32'ha8)
`define MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_1                                                         (32'hac)
`define MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_1                                                         (32'hac)
`define MCI_REG_WDT_TIMER2_EN                                                                       (32'hb0)
`define MCI_REG_WDT_TIMER2_EN                                                                       (32'hb0)
`define MCI_REG_WDT_TIMER2_EN_TIMER2_EN_LOW                                                         (0)
`define MCI_REG_WDT_TIMER2_EN_TIMER2_EN_MASK                                                        (32'h1)
`define MCI_REG_WDT_TIMER2_CTRL                                                                     (32'hb4)
`define MCI_REG_WDT_TIMER2_CTRL                                                                     (32'hb4)
`define MCI_REG_WDT_TIMER2_CTRL_TIMER2_RESTART_LOW                                                  (0)
`define MCI_REG_WDT_TIMER2_CTRL_TIMER2_RESTART_MASK                                                 (32'h1)
`define MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_0                                                         (32'hb8)
`define MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_0                                                         (32'hb8)
`define MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_1                                                         (32'hbc)
`define MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_1                                                         (32'hbc)
`define MCI_REG_WDT_STATUS                                                                          (32'hc0)
`define MCI_REG_WDT_STATUS                                                                          (32'hc0)
`define MCI_REG_WDT_STATUS_T1_TIMEOUT_LOW                                                           (0)
`define MCI_REG_WDT_STATUS_T1_TIMEOUT_MASK                                                          (32'h1)
`define MCI_REG_WDT_STATUS_T2_TIMEOUT_LOW                                                           (1)
`define MCI_REG_WDT_STATUS_T2_TIMEOUT_MASK                                                          (32'h2)
`define MCI_REG_WDT_CFG_0                                                                           (32'hd0)
`define MCI_REG_WDT_CFG_0                                                                           (32'hd0)
`define MCI_REG_WDT_CFG_1                                                                           (32'hd4)
`define MCI_REG_WDT_CFG_1                                                                           (32'hd4)
`define MCI_REG_MCU_TIMER_CONFIG                                                                    (32'he0)
`define MCI_REG_MCU_TIMER_CONFIG                                                                    (32'he0)
`define MCI_REG_MCU_RV_MTIME_L                                                                      (32'he4)
`define MCI_REG_MCU_RV_MTIME_L                                                                      (32'he4)
`define MCI_REG_MCU_RV_MTIME_H                                                                      (32'he8)
`define MCI_REG_MCU_RV_MTIME_H                                                                      (32'he8)
`define MCI_REG_MCU_RV_MTIMECMP_L                                                                   (32'hec)
`define MCI_REG_MCU_RV_MTIMECMP_L                                                                   (32'hec)
`define MCI_REG_MCU_RV_MTIMECMP_H                                                                   (32'hf0)
`define MCI_REG_MCU_RV_MTIMECMP_H                                                                   (32'hf0)
`define MCI_REG_RESET_REQUEST                                                                       (32'h100)
`define MCI_REG_RESET_REQUEST                                                                       (32'h100)
`define MCI_REG_RESET_REQUEST_MCU_REQ_LOW                                                           (0)
`define MCI_REG_RESET_REQUEST_MCU_REQ_MASK                                                          (32'h1)
`define MCI_REG_MCI_BOOTFSM_GO                                                                      (32'h104)
`define MCI_REG_MCI_BOOTFSM_GO                                                                      (32'h104)
`define MCI_REG_MCI_BOOTFSM_GO_GO_LOW                                                               (0)
`define MCI_REG_MCI_BOOTFSM_GO_GO_MASK                                                              (32'h1)
`define MCI_REG_FW_SRAM_EXEC_REGION_SIZE                                                            (32'h108)
`define MCI_REG_FW_SRAM_EXEC_REGION_SIZE                                                            (32'h108)
`define MCI_REG_FW_SRAM_EXEC_REGION_SIZE_SIZE_LOW                                                   (0)
`define MCI_REG_FW_SRAM_EXEC_REGION_SIZE_SIZE_MASK                                                  (32'hffff)
`define MCI_REG_MCU_NMI_VECTOR                                                                      (32'h10c)
`define MCI_REG_MCU_NMI_VECTOR                                                                      (32'h10c)
`define MCI_REG_MCU_RESET_VECTOR                                                                    (32'h110)
`define MCI_REG_MCU_RESET_VECTOR                                                                    (32'h110)
`define MCI_REG_MBOX0_VALID_AXI_ID_0                                                                (32'h180)
`define MCI_REG_MBOX0_VALID_AXI_ID_0                                                                (32'h180)
`define MCI_REG_MBOX0_VALID_AXI_ID_1                                                                (32'h184)
`define MCI_REG_MBOX0_VALID_AXI_ID_1                                                                (32'h184)
`define MCI_REG_MBOX0_VALID_AXI_ID_2                                                                (32'h188)
`define MCI_REG_MBOX0_VALID_AXI_ID_2                                                                (32'h188)
`define MCI_REG_MBOX0_VALID_AXI_ID_3                                                                (32'h18c)
`define MCI_REG_MBOX0_VALID_AXI_ID_3                                                                (32'h18c)
`define MCI_REG_MBOX0_VALID_AXI_ID_4                                                                (32'h190)
`define MCI_REG_MBOX0_VALID_AXI_ID_4                                                                (32'h190)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_0                                                           (32'h1a0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_0                                                           (32'h1a0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_0_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_0_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_1                                                           (32'h1a4)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_1                                                           (32'h1a4)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_1_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_1_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_2                                                           (32'h1a8)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_2                                                           (32'h1a8)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_2_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_2_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_3                                                           (32'h1ac)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_3                                                           (32'h1ac)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_3_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_3_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_4                                                           (32'h1b0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_4                                                           (32'h1b0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_4_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX0_VALID_AXI_ID_LOCK_4_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX1_VALID_AXI_ID_0                                                                (32'h1c0)
`define MCI_REG_MBOX1_VALID_AXI_ID_0                                                                (32'h1c0)
`define MCI_REG_MBOX1_VALID_AXI_ID_1                                                                (32'h1c4)
`define MCI_REG_MBOX1_VALID_AXI_ID_1                                                                (32'h1c4)
`define MCI_REG_MBOX1_VALID_AXI_ID_2                                                                (32'h1c8)
`define MCI_REG_MBOX1_VALID_AXI_ID_2                                                                (32'h1c8)
`define MCI_REG_MBOX1_VALID_AXI_ID_3                                                                (32'h1cc)
`define MCI_REG_MBOX1_VALID_AXI_ID_3                                                                (32'h1cc)
`define MCI_REG_MBOX1_VALID_AXI_ID_4                                                                (32'h1d0)
`define MCI_REG_MBOX1_VALID_AXI_ID_4                                                                (32'h1d0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_0                                                           (32'h1e0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_0                                                           (32'h1e0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_0_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_0_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_1                                                           (32'h1e4)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_1                                                           (32'h1e4)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_1_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_1_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_2                                                           (32'h1e8)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_2                                                           (32'h1e8)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_2_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_2_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_3                                                           (32'h1ec)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_3                                                           (32'h1ec)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_3_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_3_LOCK_MASK                                                 (32'h1)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_4                                                           (32'h1f0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_4                                                           (32'h1f0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_4_LOCK_LOW                                                  (0)
`define MCI_REG_MBOX1_VALID_AXI_ID_LOCK_4_LOCK_MASK                                                 (32'h1)
`define MCI_REG_GENERIC_INPUT_WIRES_0                                                               (32'h400)
`define MCI_REG_GENERIC_INPUT_WIRES_0                                                               (32'h400)
`define MCI_REG_GENERIC_INPUT_WIRES_1                                                               (32'h404)
`define MCI_REG_GENERIC_INPUT_WIRES_1                                                               (32'h404)
`define MCI_REG_GENERIC_OUTPUT_WIRES_0                                                              (32'h408)
`define MCI_REG_GENERIC_OUTPUT_WIRES_0                                                              (32'h408)
`define MCI_REG_GENERIC_OUTPUT_WIRES_1                                                              (32'h40c)
`define MCI_REG_GENERIC_OUTPUT_WIRES_1                                                              (32'h40c)
`define MCI_REG_DEBUG_IN                                                                            (32'h410)
`define MCI_REG_DEBUG_IN                                                                            (32'h410)
`define MCI_REG_DEBUG_IN_FIXME_LOW                                                                  (0)
`define MCI_REG_DEBUG_IN_FIXME_MASK                                                                 (32'h1)
`define MCI_REG_DEBUG_OUT                                                                           (32'h414)
`define MCI_REG_DEBUG_OUT                                                                           (32'h414)
`define MCI_REG_DEBUG_OUT_FIXME_LOW                                                                 (0)
`define MCI_REG_DEBUG_OUT_FIXME_MASK                                                                (32'h1)
`define MCI_REG_FUSE_WR_DONE                                                                        (32'h440)
`define MCI_REG_FUSE_WR_DONE                                                                        (32'h440)
`define MCI_REG_FUSE_WR_DONE_DONE_LOW                                                               (0)
`define MCI_REG_FUSE_WR_DONE_DONE_MASK                                                              (32'h1)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_0                                                   (32'h480)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_0                                                   (32'h480)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_1                                                   (32'h484)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_1                                                   (32'h484)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_2                                                   (32'h488)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_2                                                   (32'h488)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_3                                                   (32'h48c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_3                                                   (32'h48c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_4                                                   (32'h490)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_4                                                   (32'h490)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_5                                                   (32'h494)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_5                                                   (32'h494)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_6                                                   (32'h498)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_6                                                   (32'h498)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_7                                                   (32'h49c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_7                                                   (32'h49c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_8                                                   (32'h4a0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_8                                                   (32'h4a0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_9                                                   (32'h4a4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_9                                                   (32'h4a4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_10                                                  (32'h4a8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_10                                                  (32'h4a8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_11                                                  (32'h4ac)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_11                                                  (32'h4ac)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_0                                                   (32'h4b0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_0                                                   (32'h4b0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_1                                                   (32'h4b4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_1                                                   (32'h4b4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_2                                                   (32'h4b8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_2                                                   (32'h4b8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_3                                                   (32'h4bc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_3                                                   (32'h4bc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_4                                                   (32'h4c0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_4                                                   (32'h4c0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_5                                                   (32'h4c4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_5                                                   (32'h4c4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_6                                                   (32'h4c8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_6                                                   (32'h4c8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_7                                                   (32'h4cc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_7                                                   (32'h4cc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_8                                                   (32'h4d0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_8                                                   (32'h4d0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_9                                                   (32'h4d4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_9                                                   (32'h4d4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_10                                                  (32'h4d8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_10                                                  (32'h4d8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_11                                                  (32'h4dc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_11                                                  (32'h4dc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_0                                                   (32'h4e0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_0                                                   (32'h4e0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_1                                                   (32'h4e4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_1                                                   (32'h4e4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_2                                                   (32'h4e8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_2                                                   (32'h4e8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_3                                                   (32'h4ec)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_3                                                   (32'h4ec)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_4                                                   (32'h4f0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_4                                                   (32'h4f0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_5                                                   (32'h4f4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_5                                                   (32'h4f4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_6                                                   (32'h4f8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_6                                                   (32'h4f8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_7                                                   (32'h4fc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_7                                                   (32'h4fc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_8                                                   (32'h500)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_8                                                   (32'h500)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_9                                                   (32'h504)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_9                                                   (32'h504)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_10                                                  (32'h508)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_10                                                  (32'h508)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_11                                                  (32'h50c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_11                                                  (32'h50c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_0                                                   (32'h510)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_0                                                   (32'h510)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_1                                                   (32'h514)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_1                                                   (32'h514)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_2                                                   (32'h518)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_2                                                   (32'h518)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_3                                                   (32'h51c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_3                                                   (32'h51c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_4                                                   (32'h520)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_4                                                   (32'h520)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_5                                                   (32'h524)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_5                                                   (32'h524)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_6                                                   (32'h528)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_6                                                   (32'h528)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_7                                                   (32'h52c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_7                                                   (32'h52c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_8                                                   (32'h530)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_8                                                   (32'h530)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_9                                                   (32'h534)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_9                                                   (32'h534)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_10                                                  (32'h538)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_10                                                  (32'h538)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_11                                                  (32'h53c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_11                                                  (32'h53c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_0                                                   (32'h540)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_0                                                   (32'h540)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_1                                                   (32'h544)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_1                                                   (32'h544)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_2                                                   (32'h548)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_2                                                   (32'h548)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_3                                                   (32'h54c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_3                                                   (32'h54c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_4                                                   (32'h550)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_4                                                   (32'h550)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_5                                                   (32'h554)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_5                                                   (32'h554)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_6                                                   (32'h558)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_6                                                   (32'h558)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_7                                                   (32'h55c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_7                                                   (32'h55c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_8                                                   (32'h560)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_8                                                   (32'h560)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_9                                                   (32'h564)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_9                                                   (32'h564)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_10                                                  (32'h568)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_10                                                  (32'h568)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_11                                                  (32'h56c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_11                                                  (32'h56c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_0                                                   (32'h570)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_0                                                   (32'h570)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_1                                                   (32'h574)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_1                                                   (32'h574)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_2                                                   (32'h578)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_2                                                   (32'h578)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_3                                                   (32'h57c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_3                                                   (32'h57c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_4                                                   (32'h580)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_4                                                   (32'h580)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_5                                                   (32'h584)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_5                                                   (32'h584)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_6                                                   (32'h588)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_6                                                   (32'h588)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_7                                                   (32'h58c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_7                                                   (32'h58c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_8                                                   (32'h590)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_8                                                   (32'h590)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_9                                                   (32'h594)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_9                                                   (32'h594)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_10                                                  (32'h598)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_10                                                  (32'h598)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_11                                                  (32'h59c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_11                                                  (32'h59c)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_0                                                   (32'h5a0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_0                                                   (32'h5a0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_1                                                   (32'h5a4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_1                                                   (32'h5a4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_2                                                   (32'h5a8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_2                                                   (32'h5a8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_3                                                   (32'h5ac)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_3                                                   (32'h5ac)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_4                                                   (32'h5b0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_4                                                   (32'h5b0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_5                                                   (32'h5b4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_5                                                   (32'h5b4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_6                                                   (32'h5b8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_6                                                   (32'h5b8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_7                                                   (32'h5bc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_7                                                   (32'h5bc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_8                                                   (32'h5c0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_8                                                   (32'h5c0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_9                                                   (32'h5c4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_9                                                   (32'h5c4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_10                                                  (32'h5c8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_10                                                  (32'h5c8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_11                                                  (32'h5cc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_11                                                  (32'h5cc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_0                                                   (32'h5d0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_0                                                   (32'h5d0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_1                                                   (32'h5d4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_1                                                   (32'h5d4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_2                                                   (32'h5d8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_2                                                   (32'h5d8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_3                                                   (32'h5dc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_3                                                   (32'h5dc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_4                                                   (32'h5e0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_4                                                   (32'h5e0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_5                                                   (32'h5e4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_5                                                   (32'h5e4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_6                                                   (32'h5e8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_6                                                   (32'h5e8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_7                                                   (32'h5ec)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_7                                                   (32'h5ec)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_8                                                   (32'h5f0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_8                                                   (32'h5f0)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_9                                                   (32'h5f4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_9                                                   (32'h5f4)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_10                                                  (32'h5f8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_10                                                  (32'h5f8)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_11                                                  (32'h5fc)
`define MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_11                                                  (32'h5fc)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_0                                                            (32'h800)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_0                                                            (32'h800)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_0_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_0_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_1                                                            (32'h804)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_1                                                            (32'h804)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_1_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_1_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_2                                                            (32'h808)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_2                                                            (32'h808)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_2_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_2_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_3                                                            (32'h80c)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_3                                                            (32'h80c)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_3_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_3_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_4                                                            (32'h810)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_4                                                            (32'h810)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_4_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_4_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_5                                                            (32'h814)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_5                                                            (32'h814)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_5_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_5_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_6                                                            (32'h818)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_6                                                            (32'h818)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_6_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_6_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_7                                                            (32'h81c)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_7                                                            (32'h81c)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_7_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_7_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_8                                                            (32'h820)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_8                                                            (32'h820)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_8_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_8_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_9                                                            (32'h824)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_9                                                            (32'h824)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_9_LOCK_ENTRY_LOW                                             (0)
`define MCI_REG_STICKY_DATA_VAULT_CTRL_9_LOCK_ENTRY_MASK                                            (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                         (32'h828)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                         (32'h828)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                         (32'h82c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                         (32'h82c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                         (32'h830)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                         (32'h830)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                         (32'h834)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                         (32'h834)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                         (32'h838)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                         (32'h838)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                         (32'h83c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                         (32'h83c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                         (32'h840)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                         (32'h840)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                         (32'h844)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                         (32'h844)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                         (32'h848)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                         (32'h848)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                         (32'h84c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                         (32'h84c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                        (32'h850)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                        (32'h850)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                        (32'h854)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                        (32'h854)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_0_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                         (32'h858)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                         (32'h858)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                         (32'h85c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                         (32'h85c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                         (32'h860)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                         (32'h860)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                         (32'h864)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                         (32'h864)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                         (32'h868)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                         (32'h868)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                         (32'h86c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                         (32'h86c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                         (32'h870)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                         (32'h870)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                         (32'h874)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                         (32'h874)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                         (32'h878)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                         (32'h878)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                         (32'h87c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                         (32'h87c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                        (32'h880)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                        (32'h880)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                        (32'h884)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                        (32'h884)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_1_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                         (32'h888)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                         (32'h888)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                         (32'h88c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                         (32'h88c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                         (32'h890)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                         (32'h890)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                         (32'h894)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                         (32'h894)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                         (32'h898)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                         (32'h898)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                         (32'h89c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                         (32'h89c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                         (32'h8a0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                         (32'h8a0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                         (32'h8a4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                         (32'h8a4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                         (32'h8a8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                         (32'h8a8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                         (32'h8ac)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                         (32'h8ac)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                        (32'h8b0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                        (32'h8b0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                        (32'h8b4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                        (32'h8b4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_2_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                         (32'h8b8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                         (32'h8b8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                         (32'h8bc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                         (32'h8bc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                         (32'h8c0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                         (32'h8c0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                         (32'h8c4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                         (32'h8c4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                         (32'h8c8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                         (32'h8c8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                         (32'h8cc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                         (32'h8cc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                         (32'h8d0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                         (32'h8d0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                         (32'h8d4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                         (32'h8d4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                         (32'h8d8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                         (32'h8d8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                         (32'h8dc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                         (32'h8dc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                        (32'h8e0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                        (32'h8e0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                        (32'h8e4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                        (32'h8e4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_3_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                         (32'h8e8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                         (32'h8e8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                         (32'h8ec)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                         (32'h8ec)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                         (32'h8f0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                         (32'h8f0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                         (32'h8f4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                         (32'h8f4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                         (32'h8f8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                         (32'h8f8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                         (32'h8fc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                         (32'h8fc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                         (32'h900)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                         (32'h900)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                         (32'h904)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                         (32'h904)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                         (32'h908)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                         (32'h908)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                         (32'h90c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                         (32'h90c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                        (32'h910)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                        (32'h910)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                        (32'h914)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                        (32'h914)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_4_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                         (32'h918)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                         (32'h918)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                         (32'h91c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                         (32'h91c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                         (32'h920)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                         (32'h920)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                         (32'h924)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                         (32'h924)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                         (32'h928)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                         (32'h928)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                         (32'h92c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                         (32'h92c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                         (32'h930)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                         (32'h930)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                         (32'h934)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                         (32'h934)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                         (32'h938)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                         (32'h938)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                         (32'h93c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                         (32'h93c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                        (32'h940)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                        (32'h940)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                        (32'h944)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                        (32'h944)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_5_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                         (32'h948)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                         (32'h948)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                         (32'h94c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                         (32'h94c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                         (32'h950)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                         (32'h950)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                         (32'h954)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                         (32'h954)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                         (32'h958)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                         (32'h958)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                         (32'h95c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                         (32'h95c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                         (32'h960)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                         (32'h960)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                         (32'h964)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                         (32'h964)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                         (32'h968)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                         (32'h968)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                         (32'h96c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                         (32'h96c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                        (32'h970)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                        (32'h970)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                        (32'h974)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                        (32'h974)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_6_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                         (32'h978)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                         (32'h978)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                         (32'h97c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                         (32'h97c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                         (32'h980)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                         (32'h980)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                         (32'h984)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                         (32'h984)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                         (32'h988)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                         (32'h988)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                         (32'h98c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                         (32'h98c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                         (32'h990)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                         (32'h990)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                         (32'h994)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                         (32'h994)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                         (32'h998)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                         (32'h998)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                         (32'h99c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                         (32'h99c)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                        (32'h9a0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                        (32'h9a0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                        (32'h9a4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                        (32'h9a4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_7_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                         (32'h9a8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                         (32'h9a8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                         (32'h9ac)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                         (32'h9ac)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                         (32'h9b0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                         (32'h9b0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                         (32'h9b4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                         (32'h9b4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                         (32'h9b8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                         (32'h9b8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                         (32'h9bc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                         (32'h9bc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                         (32'h9c0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                         (32'h9c0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                         (32'h9c4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                         (32'h9c4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                         (32'h9c8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                         (32'h9c8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                         (32'h9cc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                         (32'h9cc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                        (32'h9d0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                        (32'h9d0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                        (32'h9d4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                        (32'h9d4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_8_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                         (32'h9d8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                         (32'h9d8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                         (32'h9dc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                         (32'h9dc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                         (32'h9e0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                         (32'h9e0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                         (32'h9e4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                         (32'h9e4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                         (32'h9e8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                         (32'h9e8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                         (32'h9ec)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                         (32'h9ec)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                         (32'h9f0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                         (32'h9f0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                         (32'h9f4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                         (32'h9f4)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                         (32'h9f8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                         (32'h9f8)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                         (32'h9fc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                         (32'h9fc)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                        (32'ha00)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                        (32'ha00)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_10_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_10_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                        (32'ha04)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                        (32'ha04)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_11_LOCK_ENTRY_LOW                                         (0)
`define MCI_REG_STICKY_DATA_VAULT_ENTRY_9_11_LOCK_ENTRY_MASK                                        (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_0                                                                   (32'ha08)
`define MCI_REG_DATA_VAULT_CTRL_0                                                                   (32'ha08)
`define MCI_REG_DATA_VAULT_CTRL_0_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_0_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_1                                                                   (32'ha0c)
`define MCI_REG_DATA_VAULT_CTRL_1                                                                   (32'ha0c)
`define MCI_REG_DATA_VAULT_CTRL_1_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_1_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_2                                                                   (32'ha10)
`define MCI_REG_DATA_VAULT_CTRL_2                                                                   (32'ha10)
`define MCI_REG_DATA_VAULT_CTRL_2_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_2_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_3                                                                   (32'ha14)
`define MCI_REG_DATA_VAULT_CTRL_3                                                                   (32'ha14)
`define MCI_REG_DATA_VAULT_CTRL_3_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_3_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_4                                                                   (32'ha18)
`define MCI_REG_DATA_VAULT_CTRL_4                                                                   (32'ha18)
`define MCI_REG_DATA_VAULT_CTRL_4_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_4_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_5                                                                   (32'ha1c)
`define MCI_REG_DATA_VAULT_CTRL_5                                                                   (32'ha1c)
`define MCI_REG_DATA_VAULT_CTRL_5_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_5_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_6                                                                   (32'ha20)
`define MCI_REG_DATA_VAULT_CTRL_6                                                                   (32'ha20)
`define MCI_REG_DATA_VAULT_CTRL_6_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_6_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_7                                                                   (32'ha24)
`define MCI_REG_DATA_VAULT_CTRL_7                                                                   (32'ha24)
`define MCI_REG_DATA_VAULT_CTRL_7_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_7_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_8                                                                   (32'ha28)
`define MCI_REG_DATA_VAULT_CTRL_8                                                                   (32'ha28)
`define MCI_REG_DATA_VAULT_CTRL_8_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_8_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_CTRL_9                                                                   (32'ha2c)
`define MCI_REG_DATA_VAULT_CTRL_9                                                                   (32'ha2c)
`define MCI_REG_DATA_VAULT_CTRL_9_LOCK_ENTRY_LOW                                                    (0)
`define MCI_REG_DATA_VAULT_CTRL_9_LOCK_ENTRY_MASK                                                   (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_0                                                                (32'ha30)
`define MCI_REG_DATA_VAULT_ENTRY_0_0                                                                (32'ha30)
`define MCI_REG_DATA_VAULT_ENTRY_0_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_1                                                                (32'ha34)
`define MCI_REG_DATA_VAULT_ENTRY_0_1                                                                (32'ha34)
`define MCI_REG_DATA_VAULT_ENTRY_0_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_2                                                                (32'ha38)
`define MCI_REG_DATA_VAULT_ENTRY_0_2                                                                (32'ha38)
`define MCI_REG_DATA_VAULT_ENTRY_0_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_3                                                                (32'ha3c)
`define MCI_REG_DATA_VAULT_ENTRY_0_3                                                                (32'ha3c)
`define MCI_REG_DATA_VAULT_ENTRY_0_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_4                                                                (32'ha40)
`define MCI_REG_DATA_VAULT_ENTRY_0_4                                                                (32'ha40)
`define MCI_REG_DATA_VAULT_ENTRY_0_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_5                                                                (32'ha44)
`define MCI_REG_DATA_VAULT_ENTRY_0_5                                                                (32'ha44)
`define MCI_REG_DATA_VAULT_ENTRY_0_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_6                                                                (32'ha48)
`define MCI_REG_DATA_VAULT_ENTRY_0_6                                                                (32'ha48)
`define MCI_REG_DATA_VAULT_ENTRY_0_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_7                                                                (32'ha4c)
`define MCI_REG_DATA_VAULT_ENTRY_0_7                                                                (32'ha4c)
`define MCI_REG_DATA_VAULT_ENTRY_0_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_8                                                                (32'ha50)
`define MCI_REG_DATA_VAULT_ENTRY_0_8                                                                (32'ha50)
`define MCI_REG_DATA_VAULT_ENTRY_0_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_9                                                                (32'ha54)
`define MCI_REG_DATA_VAULT_ENTRY_0_9                                                                (32'ha54)
`define MCI_REG_DATA_VAULT_ENTRY_0_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_10                                                               (32'ha58)
`define MCI_REG_DATA_VAULT_ENTRY_0_10                                                               (32'ha58)
`define MCI_REG_DATA_VAULT_ENTRY_0_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_0_11                                                               (32'ha5c)
`define MCI_REG_DATA_VAULT_ENTRY_0_11                                                               (32'ha5c)
`define MCI_REG_DATA_VAULT_ENTRY_0_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_0_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_0                                                                (32'ha60)
`define MCI_REG_DATA_VAULT_ENTRY_1_0                                                                (32'ha60)
`define MCI_REG_DATA_VAULT_ENTRY_1_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_1                                                                (32'ha64)
`define MCI_REG_DATA_VAULT_ENTRY_1_1                                                                (32'ha64)
`define MCI_REG_DATA_VAULT_ENTRY_1_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_2                                                                (32'ha68)
`define MCI_REG_DATA_VAULT_ENTRY_1_2                                                                (32'ha68)
`define MCI_REG_DATA_VAULT_ENTRY_1_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_3                                                                (32'ha6c)
`define MCI_REG_DATA_VAULT_ENTRY_1_3                                                                (32'ha6c)
`define MCI_REG_DATA_VAULT_ENTRY_1_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_4                                                                (32'ha70)
`define MCI_REG_DATA_VAULT_ENTRY_1_4                                                                (32'ha70)
`define MCI_REG_DATA_VAULT_ENTRY_1_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_5                                                                (32'ha74)
`define MCI_REG_DATA_VAULT_ENTRY_1_5                                                                (32'ha74)
`define MCI_REG_DATA_VAULT_ENTRY_1_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_6                                                                (32'ha78)
`define MCI_REG_DATA_VAULT_ENTRY_1_6                                                                (32'ha78)
`define MCI_REG_DATA_VAULT_ENTRY_1_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_7                                                                (32'ha7c)
`define MCI_REG_DATA_VAULT_ENTRY_1_7                                                                (32'ha7c)
`define MCI_REG_DATA_VAULT_ENTRY_1_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_8                                                                (32'ha80)
`define MCI_REG_DATA_VAULT_ENTRY_1_8                                                                (32'ha80)
`define MCI_REG_DATA_VAULT_ENTRY_1_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_9                                                                (32'ha84)
`define MCI_REG_DATA_VAULT_ENTRY_1_9                                                                (32'ha84)
`define MCI_REG_DATA_VAULT_ENTRY_1_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_10                                                               (32'ha88)
`define MCI_REG_DATA_VAULT_ENTRY_1_10                                                               (32'ha88)
`define MCI_REG_DATA_VAULT_ENTRY_1_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_1_11                                                               (32'ha8c)
`define MCI_REG_DATA_VAULT_ENTRY_1_11                                                               (32'ha8c)
`define MCI_REG_DATA_VAULT_ENTRY_1_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_1_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_0                                                                (32'ha90)
`define MCI_REG_DATA_VAULT_ENTRY_2_0                                                                (32'ha90)
`define MCI_REG_DATA_VAULT_ENTRY_2_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_1                                                                (32'ha94)
`define MCI_REG_DATA_VAULT_ENTRY_2_1                                                                (32'ha94)
`define MCI_REG_DATA_VAULT_ENTRY_2_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_2                                                                (32'ha98)
`define MCI_REG_DATA_VAULT_ENTRY_2_2                                                                (32'ha98)
`define MCI_REG_DATA_VAULT_ENTRY_2_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_3                                                                (32'ha9c)
`define MCI_REG_DATA_VAULT_ENTRY_2_3                                                                (32'ha9c)
`define MCI_REG_DATA_VAULT_ENTRY_2_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_4                                                                (32'haa0)
`define MCI_REG_DATA_VAULT_ENTRY_2_4                                                                (32'haa0)
`define MCI_REG_DATA_VAULT_ENTRY_2_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_5                                                                (32'haa4)
`define MCI_REG_DATA_VAULT_ENTRY_2_5                                                                (32'haa4)
`define MCI_REG_DATA_VAULT_ENTRY_2_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_6                                                                (32'haa8)
`define MCI_REG_DATA_VAULT_ENTRY_2_6                                                                (32'haa8)
`define MCI_REG_DATA_VAULT_ENTRY_2_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_7                                                                (32'haac)
`define MCI_REG_DATA_VAULT_ENTRY_2_7                                                                (32'haac)
`define MCI_REG_DATA_VAULT_ENTRY_2_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_8                                                                (32'hab0)
`define MCI_REG_DATA_VAULT_ENTRY_2_8                                                                (32'hab0)
`define MCI_REG_DATA_VAULT_ENTRY_2_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_9                                                                (32'hab4)
`define MCI_REG_DATA_VAULT_ENTRY_2_9                                                                (32'hab4)
`define MCI_REG_DATA_VAULT_ENTRY_2_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_10                                                               (32'hab8)
`define MCI_REG_DATA_VAULT_ENTRY_2_10                                                               (32'hab8)
`define MCI_REG_DATA_VAULT_ENTRY_2_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_2_11                                                               (32'habc)
`define MCI_REG_DATA_VAULT_ENTRY_2_11                                                               (32'habc)
`define MCI_REG_DATA_VAULT_ENTRY_2_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_2_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_0                                                                (32'hac0)
`define MCI_REG_DATA_VAULT_ENTRY_3_0                                                                (32'hac0)
`define MCI_REG_DATA_VAULT_ENTRY_3_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_1                                                                (32'hac4)
`define MCI_REG_DATA_VAULT_ENTRY_3_1                                                                (32'hac4)
`define MCI_REG_DATA_VAULT_ENTRY_3_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_2                                                                (32'hac8)
`define MCI_REG_DATA_VAULT_ENTRY_3_2                                                                (32'hac8)
`define MCI_REG_DATA_VAULT_ENTRY_3_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_3                                                                (32'hacc)
`define MCI_REG_DATA_VAULT_ENTRY_3_3                                                                (32'hacc)
`define MCI_REG_DATA_VAULT_ENTRY_3_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_4                                                                (32'had0)
`define MCI_REG_DATA_VAULT_ENTRY_3_4                                                                (32'had0)
`define MCI_REG_DATA_VAULT_ENTRY_3_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_5                                                                (32'had4)
`define MCI_REG_DATA_VAULT_ENTRY_3_5                                                                (32'had4)
`define MCI_REG_DATA_VAULT_ENTRY_3_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_6                                                                (32'had8)
`define MCI_REG_DATA_VAULT_ENTRY_3_6                                                                (32'had8)
`define MCI_REG_DATA_VAULT_ENTRY_3_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_7                                                                (32'hadc)
`define MCI_REG_DATA_VAULT_ENTRY_3_7                                                                (32'hadc)
`define MCI_REG_DATA_VAULT_ENTRY_3_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_8                                                                (32'hae0)
`define MCI_REG_DATA_VAULT_ENTRY_3_8                                                                (32'hae0)
`define MCI_REG_DATA_VAULT_ENTRY_3_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_9                                                                (32'hae4)
`define MCI_REG_DATA_VAULT_ENTRY_3_9                                                                (32'hae4)
`define MCI_REG_DATA_VAULT_ENTRY_3_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_10                                                               (32'hae8)
`define MCI_REG_DATA_VAULT_ENTRY_3_10                                                               (32'hae8)
`define MCI_REG_DATA_VAULT_ENTRY_3_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_3_11                                                               (32'haec)
`define MCI_REG_DATA_VAULT_ENTRY_3_11                                                               (32'haec)
`define MCI_REG_DATA_VAULT_ENTRY_3_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_3_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_0                                                                (32'haf0)
`define MCI_REG_DATA_VAULT_ENTRY_4_0                                                                (32'haf0)
`define MCI_REG_DATA_VAULT_ENTRY_4_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_1                                                                (32'haf4)
`define MCI_REG_DATA_VAULT_ENTRY_4_1                                                                (32'haf4)
`define MCI_REG_DATA_VAULT_ENTRY_4_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_2                                                                (32'haf8)
`define MCI_REG_DATA_VAULT_ENTRY_4_2                                                                (32'haf8)
`define MCI_REG_DATA_VAULT_ENTRY_4_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_3                                                                (32'hafc)
`define MCI_REG_DATA_VAULT_ENTRY_4_3                                                                (32'hafc)
`define MCI_REG_DATA_VAULT_ENTRY_4_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_4                                                                (32'hb00)
`define MCI_REG_DATA_VAULT_ENTRY_4_4                                                                (32'hb00)
`define MCI_REG_DATA_VAULT_ENTRY_4_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_5                                                                (32'hb04)
`define MCI_REG_DATA_VAULT_ENTRY_4_5                                                                (32'hb04)
`define MCI_REG_DATA_VAULT_ENTRY_4_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_6                                                                (32'hb08)
`define MCI_REG_DATA_VAULT_ENTRY_4_6                                                                (32'hb08)
`define MCI_REG_DATA_VAULT_ENTRY_4_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_7                                                                (32'hb0c)
`define MCI_REG_DATA_VAULT_ENTRY_4_7                                                                (32'hb0c)
`define MCI_REG_DATA_VAULT_ENTRY_4_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_8                                                                (32'hb10)
`define MCI_REG_DATA_VAULT_ENTRY_4_8                                                                (32'hb10)
`define MCI_REG_DATA_VAULT_ENTRY_4_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_9                                                                (32'hb14)
`define MCI_REG_DATA_VAULT_ENTRY_4_9                                                                (32'hb14)
`define MCI_REG_DATA_VAULT_ENTRY_4_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_10                                                               (32'hb18)
`define MCI_REG_DATA_VAULT_ENTRY_4_10                                                               (32'hb18)
`define MCI_REG_DATA_VAULT_ENTRY_4_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_4_11                                                               (32'hb1c)
`define MCI_REG_DATA_VAULT_ENTRY_4_11                                                               (32'hb1c)
`define MCI_REG_DATA_VAULT_ENTRY_4_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_4_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_0                                                                (32'hb20)
`define MCI_REG_DATA_VAULT_ENTRY_5_0                                                                (32'hb20)
`define MCI_REG_DATA_VAULT_ENTRY_5_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_1                                                                (32'hb24)
`define MCI_REG_DATA_VAULT_ENTRY_5_1                                                                (32'hb24)
`define MCI_REG_DATA_VAULT_ENTRY_5_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_2                                                                (32'hb28)
`define MCI_REG_DATA_VAULT_ENTRY_5_2                                                                (32'hb28)
`define MCI_REG_DATA_VAULT_ENTRY_5_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_3                                                                (32'hb2c)
`define MCI_REG_DATA_VAULT_ENTRY_5_3                                                                (32'hb2c)
`define MCI_REG_DATA_VAULT_ENTRY_5_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_4                                                                (32'hb30)
`define MCI_REG_DATA_VAULT_ENTRY_5_4                                                                (32'hb30)
`define MCI_REG_DATA_VAULT_ENTRY_5_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_5                                                                (32'hb34)
`define MCI_REG_DATA_VAULT_ENTRY_5_5                                                                (32'hb34)
`define MCI_REG_DATA_VAULT_ENTRY_5_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_6                                                                (32'hb38)
`define MCI_REG_DATA_VAULT_ENTRY_5_6                                                                (32'hb38)
`define MCI_REG_DATA_VAULT_ENTRY_5_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_7                                                                (32'hb3c)
`define MCI_REG_DATA_VAULT_ENTRY_5_7                                                                (32'hb3c)
`define MCI_REG_DATA_VAULT_ENTRY_5_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_8                                                                (32'hb40)
`define MCI_REG_DATA_VAULT_ENTRY_5_8                                                                (32'hb40)
`define MCI_REG_DATA_VAULT_ENTRY_5_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_9                                                                (32'hb44)
`define MCI_REG_DATA_VAULT_ENTRY_5_9                                                                (32'hb44)
`define MCI_REG_DATA_VAULT_ENTRY_5_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_10                                                               (32'hb48)
`define MCI_REG_DATA_VAULT_ENTRY_5_10                                                               (32'hb48)
`define MCI_REG_DATA_VAULT_ENTRY_5_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_5_11                                                               (32'hb4c)
`define MCI_REG_DATA_VAULT_ENTRY_5_11                                                               (32'hb4c)
`define MCI_REG_DATA_VAULT_ENTRY_5_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_5_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_0                                                                (32'hb50)
`define MCI_REG_DATA_VAULT_ENTRY_6_0                                                                (32'hb50)
`define MCI_REG_DATA_VAULT_ENTRY_6_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_1                                                                (32'hb54)
`define MCI_REG_DATA_VAULT_ENTRY_6_1                                                                (32'hb54)
`define MCI_REG_DATA_VAULT_ENTRY_6_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_2                                                                (32'hb58)
`define MCI_REG_DATA_VAULT_ENTRY_6_2                                                                (32'hb58)
`define MCI_REG_DATA_VAULT_ENTRY_6_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_3                                                                (32'hb5c)
`define MCI_REG_DATA_VAULT_ENTRY_6_3                                                                (32'hb5c)
`define MCI_REG_DATA_VAULT_ENTRY_6_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_4                                                                (32'hb60)
`define MCI_REG_DATA_VAULT_ENTRY_6_4                                                                (32'hb60)
`define MCI_REG_DATA_VAULT_ENTRY_6_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_5                                                                (32'hb64)
`define MCI_REG_DATA_VAULT_ENTRY_6_5                                                                (32'hb64)
`define MCI_REG_DATA_VAULT_ENTRY_6_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_6                                                                (32'hb68)
`define MCI_REG_DATA_VAULT_ENTRY_6_6                                                                (32'hb68)
`define MCI_REG_DATA_VAULT_ENTRY_6_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_7                                                                (32'hb6c)
`define MCI_REG_DATA_VAULT_ENTRY_6_7                                                                (32'hb6c)
`define MCI_REG_DATA_VAULT_ENTRY_6_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_8                                                                (32'hb70)
`define MCI_REG_DATA_VAULT_ENTRY_6_8                                                                (32'hb70)
`define MCI_REG_DATA_VAULT_ENTRY_6_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_9                                                                (32'hb74)
`define MCI_REG_DATA_VAULT_ENTRY_6_9                                                                (32'hb74)
`define MCI_REG_DATA_VAULT_ENTRY_6_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_10                                                               (32'hb78)
`define MCI_REG_DATA_VAULT_ENTRY_6_10                                                               (32'hb78)
`define MCI_REG_DATA_VAULT_ENTRY_6_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_6_11                                                               (32'hb7c)
`define MCI_REG_DATA_VAULT_ENTRY_6_11                                                               (32'hb7c)
`define MCI_REG_DATA_VAULT_ENTRY_6_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_6_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_0                                                                (32'hb80)
`define MCI_REG_DATA_VAULT_ENTRY_7_0                                                                (32'hb80)
`define MCI_REG_DATA_VAULT_ENTRY_7_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_1                                                                (32'hb84)
`define MCI_REG_DATA_VAULT_ENTRY_7_1                                                                (32'hb84)
`define MCI_REG_DATA_VAULT_ENTRY_7_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_2                                                                (32'hb88)
`define MCI_REG_DATA_VAULT_ENTRY_7_2                                                                (32'hb88)
`define MCI_REG_DATA_VAULT_ENTRY_7_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_3                                                                (32'hb8c)
`define MCI_REG_DATA_VAULT_ENTRY_7_3                                                                (32'hb8c)
`define MCI_REG_DATA_VAULT_ENTRY_7_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_4                                                                (32'hb90)
`define MCI_REG_DATA_VAULT_ENTRY_7_4                                                                (32'hb90)
`define MCI_REG_DATA_VAULT_ENTRY_7_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_5                                                                (32'hb94)
`define MCI_REG_DATA_VAULT_ENTRY_7_5                                                                (32'hb94)
`define MCI_REG_DATA_VAULT_ENTRY_7_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_6                                                                (32'hb98)
`define MCI_REG_DATA_VAULT_ENTRY_7_6                                                                (32'hb98)
`define MCI_REG_DATA_VAULT_ENTRY_7_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_7                                                                (32'hb9c)
`define MCI_REG_DATA_VAULT_ENTRY_7_7                                                                (32'hb9c)
`define MCI_REG_DATA_VAULT_ENTRY_7_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_8                                                                (32'hba0)
`define MCI_REG_DATA_VAULT_ENTRY_7_8                                                                (32'hba0)
`define MCI_REG_DATA_VAULT_ENTRY_7_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_9                                                                (32'hba4)
`define MCI_REG_DATA_VAULT_ENTRY_7_9                                                                (32'hba4)
`define MCI_REG_DATA_VAULT_ENTRY_7_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_10                                                               (32'hba8)
`define MCI_REG_DATA_VAULT_ENTRY_7_10                                                               (32'hba8)
`define MCI_REG_DATA_VAULT_ENTRY_7_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_7_11                                                               (32'hbac)
`define MCI_REG_DATA_VAULT_ENTRY_7_11                                                               (32'hbac)
`define MCI_REG_DATA_VAULT_ENTRY_7_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_7_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_0                                                                (32'hbb0)
`define MCI_REG_DATA_VAULT_ENTRY_8_0                                                                (32'hbb0)
`define MCI_REG_DATA_VAULT_ENTRY_8_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_1                                                                (32'hbb4)
`define MCI_REG_DATA_VAULT_ENTRY_8_1                                                                (32'hbb4)
`define MCI_REG_DATA_VAULT_ENTRY_8_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_2                                                                (32'hbb8)
`define MCI_REG_DATA_VAULT_ENTRY_8_2                                                                (32'hbb8)
`define MCI_REG_DATA_VAULT_ENTRY_8_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_3                                                                (32'hbbc)
`define MCI_REG_DATA_VAULT_ENTRY_8_3                                                                (32'hbbc)
`define MCI_REG_DATA_VAULT_ENTRY_8_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_4                                                                (32'hbc0)
`define MCI_REG_DATA_VAULT_ENTRY_8_4                                                                (32'hbc0)
`define MCI_REG_DATA_VAULT_ENTRY_8_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_5                                                                (32'hbc4)
`define MCI_REG_DATA_VAULT_ENTRY_8_5                                                                (32'hbc4)
`define MCI_REG_DATA_VAULT_ENTRY_8_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_6                                                                (32'hbc8)
`define MCI_REG_DATA_VAULT_ENTRY_8_6                                                                (32'hbc8)
`define MCI_REG_DATA_VAULT_ENTRY_8_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_7                                                                (32'hbcc)
`define MCI_REG_DATA_VAULT_ENTRY_8_7                                                                (32'hbcc)
`define MCI_REG_DATA_VAULT_ENTRY_8_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_8                                                                (32'hbd0)
`define MCI_REG_DATA_VAULT_ENTRY_8_8                                                                (32'hbd0)
`define MCI_REG_DATA_VAULT_ENTRY_8_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_9                                                                (32'hbd4)
`define MCI_REG_DATA_VAULT_ENTRY_8_9                                                                (32'hbd4)
`define MCI_REG_DATA_VAULT_ENTRY_8_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_10                                                               (32'hbd8)
`define MCI_REG_DATA_VAULT_ENTRY_8_10                                                               (32'hbd8)
`define MCI_REG_DATA_VAULT_ENTRY_8_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_8_11                                                               (32'hbdc)
`define MCI_REG_DATA_VAULT_ENTRY_8_11                                                               (32'hbdc)
`define MCI_REG_DATA_VAULT_ENTRY_8_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_8_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_0                                                                (32'hbe0)
`define MCI_REG_DATA_VAULT_ENTRY_9_0                                                                (32'hbe0)
`define MCI_REG_DATA_VAULT_ENTRY_9_0_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_0_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_1                                                                (32'hbe4)
`define MCI_REG_DATA_VAULT_ENTRY_9_1                                                                (32'hbe4)
`define MCI_REG_DATA_VAULT_ENTRY_9_1_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_1_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_2                                                                (32'hbe8)
`define MCI_REG_DATA_VAULT_ENTRY_9_2                                                                (32'hbe8)
`define MCI_REG_DATA_VAULT_ENTRY_9_2_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_2_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_3                                                                (32'hbec)
`define MCI_REG_DATA_VAULT_ENTRY_9_3                                                                (32'hbec)
`define MCI_REG_DATA_VAULT_ENTRY_9_3_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_3_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_4                                                                (32'hbf0)
`define MCI_REG_DATA_VAULT_ENTRY_9_4                                                                (32'hbf0)
`define MCI_REG_DATA_VAULT_ENTRY_9_4_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_4_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_5                                                                (32'hbf4)
`define MCI_REG_DATA_VAULT_ENTRY_9_5                                                                (32'hbf4)
`define MCI_REG_DATA_VAULT_ENTRY_9_5_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_5_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_6                                                                (32'hbf8)
`define MCI_REG_DATA_VAULT_ENTRY_9_6                                                                (32'hbf8)
`define MCI_REG_DATA_VAULT_ENTRY_9_6_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_6_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_7                                                                (32'hbfc)
`define MCI_REG_DATA_VAULT_ENTRY_9_7                                                                (32'hbfc)
`define MCI_REG_DATA_VAULT_ENTRY_9_7_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_7_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_8                                                                (32'hc00)
`define MCI_REG_DATA_VAULT_ENTRY_9_8                                                                (32'hc00)
`define MCI_REG_DATA_VAULT_ENTRY_9_8_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_8_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_9                                                                (32'hc04)
`define MCI_REG_DATA_VAULT_ENTRY_9_9                                                                (32'hc04)
`define MCI_REG_DATA_VAULT_ENTRY_9_9_LOCK_ENTRY_LOW                                                 (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_9_LOCK_ENTRY_MASK                                                (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_10                                                               (32'hc08)
`define MCI_REG_DATA_VAULT_ENTRY_9_10                                                               (32'hc08)
`define MCI_REG_DATA_VAULT_ENTRY_9_10_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_10_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_DATA_VAULT_ENTRY_9_11                                                               (32'hc0c)
`define MCI_REG_DATA_VAULT_ENTRY_9_11                                                               (32'hc0c)
`define MCI_REG_DATA_VAULT_ENTRY_9_11_LOCK_ENTRY_LOW                                                (0)
`define MCI_REG_DATA_VAULT_ENTRY_9_11_LOCK_ENTRY_MASK                                               (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_0                                                  (32'hc10)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_0                                                  (32'hc10)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_0_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_0_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_1                                                  (32'hc14)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_1                                                  (32'hc14)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_1_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_1_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_2                                                  (32'hc18)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_2                                                  (32'hc18)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_2_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_2_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_3                                                  (32'hc1c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_3                                                  (32'hc1c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_3_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_3_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_4                                                  (32'hc20)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_4                                                  (32'hc20)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_4_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_4_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_5                                                  (32'hc24)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_5                                                  (32'hc24)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_5_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_5_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_6                                                  (32'hc28)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_6                                                  (32'hc28)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_6_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_6_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_7                                                  (32'hc2c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_7                                                  (32'hc2c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_7_LOCK_ENTRY_LOW                                   (0)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_CTRL_7_LOCK_ENTRY_MASK                                  (32'h1)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_0                                                       (32'hc30)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_0                                                       (32'hc30)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_1                                                       (32'hc34)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_1                                                       (32'hc34)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_2                                                       (32'hc38)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_2                                                       (32'hc38)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_3                                                       (32'hc3c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_3                                                       (32'hc3c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_4                                                       (32'hc40)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_4                                                       (32'hc40)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_5                                                       (32'hc44)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_5                                                       (32'hc44)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_6                                                       (32'hc48)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_6                                                       (32'hc48)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_7                                                       (32'hc4c)
`define MCI_REG_STICKY_LOCKABLE_SCRATCH_REG_7                                                       (32'hc4c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_0                                                         (32'hc50)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_0                                                         (32'hc50)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_0_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_0_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_1                                                         (32'hc54)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_1                                                         (32'hc54)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_1_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_1_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_2                                                         (32'hc58)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_2                                                         (32'hc58)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_2_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_2_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_3                                                         (32'hc5c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_3                                                         (32'hc5c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_3_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_3_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_4                                                         (32'hc60)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_4                                                         (32'hc60)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_4_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_4_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_5                                                         (32'hc64)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_5                                                         (32'hc64)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_5_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_5_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_6                                                         (32'hc68)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_6                                                         (32'hc68)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_6_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_6_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_7                                                         (32'hc6c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_7                                                         (32'hc6c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_7_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_7_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_8                                                         (32'hc70)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_8                                                         (32'hc70)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_8_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_8_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_9                                                         (32'hc74)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_9                                                         (32'hc74)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_9_LOCK_ENTRY_LOW                                          (0)
`define MCI_REG_LOCKABLE_SCRATCH_REG_CTRL_9_LOCK_ENTRY_MASK                                         (32'h1)
`define MCI_REG_LOCKABLE_SCRATCH_REG_0                                                              (32'hc78)
`define MCI_REG_LOCKABLE_SCRATCH_REG_0                                                              (32'hc78)
`define MCI_REG_LOCKABLE_SCRATCH_REG_1                                                              (32'hc7c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_1                                                              (32'hc7c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_2                                                              (32'hc80)
`define MCI_REG_LOCKABLE_SCRATCH_REG_2                                                              (32'hc80)
`define MCI_REG_LOCKABLE_SCRATCH_REG_3                                                              (32'hc84)
`define MCI_REG_LOCKABLE_SCRATCH_REG_3                                                              (32'hc84)
`define MCI_REG_LOCKABLE_SCRATCH_REG_4                                                              (32'hc88)
`define MCI_REG_LOCKABLE_SCRATCH_REG_4                                                              (32'hc88)
`define MCI_REG_LOCKABLE_SCRATCH_REG_5                                                              (32'hc8c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_5                                                              (32'hc8c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_6                                                              (32'hc90)
`define MCI_REG_LOCKABLE_SCRATCH_REG_6                                                              (32'hc90)
`define MCI_REG_LOCKABLE_SCRATCH_REG_7                                                              (32'hc94)
`define MCI_REG_LOCKABLE_SCRATCH_REG_7                                                              (32'hc94)
`define MCI_REG_LOCKABLE_SCRATCH_REG_8                                                              (32'hc98)
`define MCI_REG_LOCKABLE_SCRATCH_REG_8                                                              (32'hc98)
`define MCI_REG_LOCKABLE_SCRATCH_REG_9                                                              (32'hc9c)
`define MCI_REG_LOCKABLE_SCRATCH_REG_9                                                              (32'hc9c)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_0                                                    (32'hca0)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_0                                                    (32'hca0)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_1                                                    (32'hca4)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_1                                                    (32'hca4)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_2                                                    (32'hca8)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_2                                                    (32'hca8)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_3                                                    (32'hcac)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_3                                                    (32'hcac)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_4                                                    (32'hcb0)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_4                                                    (32'hcb0)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_5                                                    (32'hcb4)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_5                                                    (32'hcb4)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_6                                                    (32'hcb8)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_6                                                    (32'hcb8)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_7                                                    (32'hcbc)
`define MCI_REG_NON_STICKY_GENERIC_SCRATCH_REG_7                                                    (32'hcbc)
`define MCI_REG_INTR_BLOCK_RF_START                                                                 (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R                                                      (32'h1004)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R                                                      (32'h1004)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R_ERROR_WDT_TIMER1_TIMEOUT_EN_LOW                      (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R_ERROR_WDT_TIMER1_TIMEOUT_EN_MASK                     (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R_ERROR_WDT_TIMER2_TIMEOUT_EN_LOW                      (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R_ERROR_WDT_TIMER2_TIMEOUT_EN_MASK                     (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R                                                      (32'h1008)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R                                                      (32'h1008)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL31_EN_LOW                       (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL31_EN_MASK                      (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL30_EN_LOW                       (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL30_EN_MASK                      (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL29_EN_LOW                       (2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL29_EN_MASK                      (32'h4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL28_EN_LOW                       (3)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL28_EN_MASK                      (32'h8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL27_EN_LOW                       (4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL27_EN_MASK                      (32'h10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL26_EN_LOW                       (5)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL26_EN_MASK                      (32'h20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL25_EN_LOW                       (6)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL25_EN_MASK                      (32'h40)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL24_EN_LOW                       (7)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL24_EN_MASK                      (32'h80)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL23_EN_LOW                       (8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL23_EN_MASK                      (32'h100)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL22_EN_LOW                       (9)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL22_EN_MASK                      (32'h200)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL21_EN_LOW                       (10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL21_EN_MASK                      (32'h400)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL20_EN_LOW                       (11)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL20_EN_MASK                      (32'h800)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL19_EN_LOW                       (12)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL19_EN_MASK                      (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL18_EN_LOW                       (13)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL18_EN_MASK                      (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL17_EN_LOW                       (14)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL17_EN_MASK                      (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL16_EN_LOW                       (15)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL16_EN_MASK                      (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL15_EN_LOW                       (16)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL15_EN_MASK                      (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL14_EN_LOW                       (17)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL14_EN_MASK                      (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL13_EN_LOW                       (18)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL13_EN_MASK                      (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL12_EN_LOW                       (19)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL12_EN_MASK                      (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL11_EN_LOW                       (20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL11_EN_MASK                      (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL10_EN_LOW                       (21)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL10_EN_MASK                      (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL9_EN_LOW                        (22)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL9_EN_MASK                       (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL8_EN_LOW                        (23)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL8_EN_MASK                       (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL7_EN_LOW                        (24)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL7_EN_MASK                       (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL6_EN_LOW                        (25)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL6_EN_MASK                       (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL5_EN_LOW                        (26)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL5_EN_MASK                       (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL4_EN_LOW                        (27)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL4_EN_MASK                       (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL3_EN_LOW                        (28)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL3_EN_MASK                       (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL2_EN_LOW                        (29)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL2_EN_MASK                       (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL1_EN_LOW                        (30)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL1_EN_MASK                       (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL0_EN_LOW                        (31)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R_ERROR_AGG_ERROR_FATAL0_EN_MASK                       (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R                                                      (32'h100c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R                                                      (32'h100c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R_NOTIF_MCU_SRAM_ECC_COR_EN_LOW                        (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R_NOTIF_MCU_SRAM_ECC_COR_EN_MASK                       (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R_NOTIF_CLPRA_MCU_RESET_REQ_EN_LOW                     (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R_NOTIF_CLPRA_MCU_RESET_REQ_EN_MASK                    (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R                                                      (32'h1010)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R                                                      (32'h1010)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL31_EN_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL31_EN_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL30_EN_LOW                   (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL30_EN_MASK                  (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL29_EN_LOW                   (2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL29_EN_MASK                  (32'h4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL28_EN_LOW                   (3)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL28_EN_MASK                  (32'h8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL27_EN_LOW                   (4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL27_EN_MASK                  (32'h10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL26_EN_LOW                   (5)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL26_EN_MASK                  (32'h20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL25_EN_LOW                   (6)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL25_EN_MASK                  (32'h40)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL24_EN_LOW                   (7)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL24_EN_MASK                  (32'h80)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL23_EN_LOW                   (8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL23_EN_MASK                  (32'h100)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL22_EN_LOW                   (9)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL22_EN_MASK                  (32'h200)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL21_EN_LOW                   (10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL21_EN_MASK                  (32'h400)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL20_EN_LOW                   (11)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL20_EN_MASK                  (32'h800)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL19_EN_LOW                   (12)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL19_EN_MASK                  (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL18_EN_LOW                   (13)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL18_EN_MASK                  (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL17_EN_LOW                   (14)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL17_EN_MASK                  (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL16_EN_LOW                   (15)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL16_EN_MASK                  (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL15_EN_LOW                   (16)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL15_EN_MASK                  (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL14_EN_LOW                   (17)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL14_EN_MASK                  (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL13_EN_LOW                   (18)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL13_EN_MASK                  (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL12_EN_LOW                   (19)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL12_EN_MASK                  (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL11_EN_LOW                   (20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL11_EN_MASK                  (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL10_EN_LOW                   (21)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL10_EN_MASK                  (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL9_EN_LOW                    (22)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL9_EN_MASK                   (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL8_EN_LOW                    (23)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL8_EN_MASK                   (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL7_EN_LOW                    (24)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL7_EN_MASK                   (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL6_EN_LOW                    (25)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL6_EN_MASK                   (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL5_EN_LOW                    (26)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL5_EN_MASK                   (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL4_EN_LOW                    (27)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL4_EN_MASK                   (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL3_EN_LOW                    (28)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL3_EN_MASK                   (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL2_EN_LOW                    (29)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL2_EN_MASK                   (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL1_EN_LOW                    (30)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL1_EN_MASK                   (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL0_EN_LOW                    (31)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R_NOTIF_AGG_ERROR_NON_FATAL0_EN_MASK                   (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h1014)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h1014)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS0_LOW                                      (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS0_MASK                                     (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS1_LOW                                      (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS1_MASK                                     (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h1018)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h1018)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS0_LOW                                      (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS0_MASK                                     (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS1_LOW                                      (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS1_MASK                                     (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R                                                (32'h101c)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R                                                (32'h101c)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R_ERROR_WDT_TIMER1_TIMEOUT_STS_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R_ERROR_WDT_TIMER1_TIMEOUT_STS_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R_ERROR_WDT_TIMER2_TIMEOUT_STS_LOW               (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R_ERROR_WDT_TIMER2_TIMEOUT_STS_MASK              (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R                                                (32'h1020)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R                                                (32'h1020)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL31_STS_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL31_STS_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL30_STS_LOW                (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL30_STS_MASK               (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL29_STS_LOW                (2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL29_STS_MASK               (32'h4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL28_STS_LOW                (3)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL28_STS_MASK               (32'h8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL27_STS_LOW                (4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL27_STS_MASK               (32'h10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL26_STS_LOW                (5)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL26_STS_MASK               (32'h20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL25_STS_LOW                (6)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL25_STS_MASK               (32'h40)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL24_STS_LOW                (7)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL24_STS_MASK               (32'h80)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL23_STS_LOW                (8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL23_STS_MASK               (32'h100)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL22_STS_LOW                (9)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL22_STS_MASK               (32'h200)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL21_STS_LOW                (10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL21_STS_MASK               (32'h400)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL20_STS_LOW                (11)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL20_STS_MASK               (32'h800)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL19_STS_LOW                (12)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL19_STS_MASK               (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL18_STS_LOW                (13)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL18_STS_MASK               (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL17_STS_LOW                (14)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL17_STS_MASK               (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL16_STS_LOW                (15)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL16_STS_MASK               (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL15_STS_LOW                (16)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL15_STS_MASK               (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL14_STS_LOW                (17)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL14_STS_MASK               (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL13_STS_LOW                (18)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL13_STS_MASK               (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL12_STS_LOW                (19)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL12_STS_MASK               (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL11_STS_LOW                (20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL11_STS_MASK               (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL10_STS_LOW                (21)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL10_STS_MASK               (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL9_STS_LOW                 (22)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL9_STS_MASK                (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL8_STS_LOW                 (23)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL8_STS_MASK                (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL7_STS_LOW                 (24)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL7_STS_MASK                (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL6_STS_LOW                 (25)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL6_STS_MASK                (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL5_STS_LOW                 (26)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL5_STS_MASK                (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL4_STS_LOW                 (27)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL4_STS_MASK                (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL3_STS_LOW                 (28)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL3_STS_MASK                (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL2_STS_LOW                 (29)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL2_STS_MASK                (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL1_STS_LOW                 (30)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL1_STS_MASK                (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL0_STS_LOW                 (31)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R_ERROR_AGG_ERROR_FATAL0_STS_MASK                (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R                                                (32'h1024)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R                                                (32'h1024)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R_NOTIF_MCU_SRAM_ECC_COR_STS_LOW                 (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R_NOTIF_MCU_SRAM_ECC_COR_STS_MASK                (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R_NOTIF_CLPRA_MCU_RESET_REQ_STS_LOW              (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R_NOTIF_CLPRA_MCU_RESET_REQ_STS_MASK             (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R                                                (32'h1028)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R                                                (32'h1028)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL31_STS_LOW            (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL31_STS_MASK           (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL30_STS_LOW            (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL30_STS_MASK           (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL29_STS_LOW            (2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL29_STS_MASK           (32'h4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL28_STS_LOW            (3)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL28_STS_MASK           (32'h8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL27_STS_LOW            (4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL27_STS_MASK           (32'h10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL26_STS_LOW            (5)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL26_STS_MASK           (32'h20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL25_STS_LOW            (6)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL25_STS_MASK           (32'h40)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL24_STS_LOW            (7)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL24_STS_MASK           (32'h80)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL23_STS_LOW            (8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL23_STS_MASK           (32'h100)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL22_STS_LOW            (9)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL22_STS_MASK           (32'h200)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL21_STS_LOW            (10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL21_STS_MASK           (32'h400)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL20_STS_LOW            (11)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL20_STS_MASK           (32'h800)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL19_STS_LOW            (12)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL19_STS_MASK           (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL18_STS_LOW            (13)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL18_STS_MASK           (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL17_STS_LOW            (14)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL17_STS_MASK           (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL16_STS_LOW            (15)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL16_STS_MASK           (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL15_STS_LOW            (16)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL15_STS_MASK           (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL14_STS_LOW            (17)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL14_STS_MASK           (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL13_STS_LOW            (18)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL13_STS_MASK           (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL12_STS_LOW            (19)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL12_STS_MASK           (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL11_STS_LOW            (20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL11_STS_MASK           (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL10_STS_LOW            (21)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL10_STS_MASK           (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL9_STS_LOW             (22)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL9_STS_MASK            (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL8_STS_LOW             (23)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL8_STS_MASK            (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL7_STS_LOW             (24)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL7_STS_MASK            (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL6_STS_LOW             (25)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL6_STS_MASK            (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL5_STS_LOW             (26)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL5_STS_MASK            (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL4_STS_LOW             (27)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL4_STS_MASK            (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL3_STS_LOW             (28)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL3_STS_MASK            (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL2_STS_LOW             (29)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL2_STS_MASK            (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL1_STS_LOW             (30)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL1_STS_MASK            (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL0_STS_LOW             (31)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R_NOTIF_AGG_ERROR_NON_FATAL0_STS_MASK            (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R                                                    (32'h102c)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R                                                    (32'h102c)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R_ERROR_WDT_TIMER1_TIMEOUT_TRIG_LOW                  (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R_ERROR_WDT_TIMER1_TIMEOUT_TRIG_MASK                 (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R_ERROR_WDT_TIMER2_TIMEOUT_TRIG_LOW                  (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R_ERROR_WDT_TIMER2_TIMEOUT_TRIG_MASK                 (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R                                                    (32'h1030)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R                                                    (32'h1030)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL31_TRIG_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL31_TRIG_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL30_TRIG_LOW                   (1)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL30_TRIG_MASK                  (32'h2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL29_TRIG_LOW                   (2)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL29_TRIG_MASK                  (32'h4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL28_TRIG_LOW                   (3)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL28_TRIG_MASK                  (32'h8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL27_TRIG_LOW                   (4)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL27_TRIG_MASK                  (32'h10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL26_TRIG_LOW                   (5)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL26_TRIG_MASK                  (32'h20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL25_TRIG_LOW                   (6)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL25_TRIG_MASK                  (32'h40)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL24_TRIG_LOW                   (7)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL24_TRIG_MASK                  (32'h80)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL23_TRIG_LOW                   (8)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL23_TRIG_MASK                  (32'h100)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL22_TRIG_LOW                   (9)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL22_TRIG_MASK                  (32'h200)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL21_TRIG_LOW                   (10)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL21_TRIG_MASK                  (32'h400)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL20_TRIG_LOW                   (11)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL20_TRIG_MASK                  (32'h800)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL19_TRIG_LOW                   (12)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL19_TRIG_MASK                  (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL18_TRIG_LOW                   (13)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL18_TRIG_MASK                  (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL17_TRIG_LOW                   (14)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL17_TRIG_MASK                  (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL16_TRIG_LOW                   (15)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL16_TRIG_MASK                  (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL15_TRIG_LOW                   (16)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL15_TRIG_MASK                  (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL14_TRIG_LOW                   (17)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL14_TRIG_MASK                  (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL13_TRIG_LOW                   (18)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL13_TRIG_MASK                  (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL12_TRIG_LOW                   (19)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL12_TRIG_MASK                  (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL11_TRIG_LOW                   (20)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL11_TRIG_MASK                  (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL10_TRIG_LOW                   (21)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL10_TRIG_MASK                  (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL9_TRIG_LOW                    (22)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL9_TRIG_MASK                   (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL8_TRIG_LOW                    (23)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL8_TRIG_MASK                   (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL7_TRIG_LOW                    (24)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL7_TRIG_MASK                   (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL6_TRIG_LOW                    (25)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL6_TRIG_MASK                   (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL5_TRIG_LOW                    (26)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL5_TRIG_MASK                   (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL4_TRIG_LOW                    (27)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL4_TRIG_MASK                   (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL3_TRIG_LOW                    (28)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL3_TRIG_MASK                   (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL2_TRIG_LOW                    (29)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL2_TRIG_MASK                   (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL1_TRIG_LOW                    (30)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL1_TRIG_MASK                   (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL0_TRIG_LOW                    (31)
`define MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R_ERROR_AGG_ERROR_FATAL0_TRIG_MASK                   (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R                                                    (32'h1034)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R                                                    (32'h1034)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R_NOTIF_MCU_SRAM_ECC_COR_TRIG_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R_NOTIF_MCU_SRAM_ECC_COR_TRIG_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R_NOTIF_CLPRA_MCU_RESET_REQ_TRIG_LOW                 (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R_NOTIF_CLPRA_MCU_RESET_REQ_TRIG_MASK                (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R                                                    (32'h1038)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R                                                    (32'h1038)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL31_TRIG_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL31_TRIG_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL30_TRIG_LOW               (1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL30_TRIG_MASK              (32'h2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL29_TRIG_LOW               (2)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL29_TRIG_MASK              (32'h4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL28_TRIG_LOW               (3)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL28_TRIG_MASK              (32'h8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL27_TRIG_LOW               (4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL27_TRIG_MASK              (32'h10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL26_TRIG_LOW               (5)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL26_TRIG_MASK              (32'h20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL25_TRIG_LOW               (6)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL25_TRIG_MASK              (32'h40)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL24_TRIG_LOW               (7)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL24_TRIG_MASK              (32'h80)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL23_TRIG_LOW               (8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL23_TRIG_MASK              (32'h100)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL22_TRIG_LOW               (9)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL22_TRIG_MASK              (32'h200)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL21_TRIG_LOW               (10)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL21_TRIG_MASK              (32'h400)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL20_TRIG_LOW               (11)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL20_TRIG_MASK              (32'h800)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL19_TRIG_LOW               (12)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL19_TRIG_MASK              (32'h1000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL18_TRIG_LOW               (13)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL18_TRIG_MASK              (32'h2000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL17_TRIG_LOW               (14)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL17_TRIG_MASK              (32'h4000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL16_TRIG_LOW               (15)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL16_TRIG_MASK              (32'h8000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL15_TRIG_LOW               (16)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL15_TRIG_MASK              (32'h10000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL14_TRIG_LOW               (17)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL14_TRIG_MASK              (32'h20000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL13_TRIG_LOW               (18)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL13_TRIG_MASK              (32'h40000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL12_TRIG_LOW               (19)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL12_TRIG_MASK              (32'h80000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL11_TRIG_LOW               (20)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL11_TRIG_MASK              (32'h100000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL10_TRIG_LOW               (21)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL10_TRIG_MASK              (32'h200000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL9_TRIG_LOW                (22)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL9_TRIG_MASK               (32'h400000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL8_TRIG_LOW                (23)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL8_TRIG_MASK               (32'h800000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL7_TRIG_LOW                (24)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL7_TRIG_MASK               (32'h1000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL6_TRIG_LOW                (25)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL6_TRIG_MASK               (32'h2000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL5_TRIG_LOW                (26)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL5_TRIG_MASK               (32'h4000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL4_TRIG_LOW                (27)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL4_TRIG_MASK               (32'h8000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL3_TRIG_LOW                (28)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL3_TRIG_MASK               (32'h10000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL2_TRIG_LOW                (29)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL2_TRIG_MASK               (32'h20000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL1_TRIG_LOW                (30)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL1_TRIG_MASK               (32'h40000000)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL0_TRIG_LOW                (31)
`define MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R_NOTIF_AGG_ERROR_NON_FATAL0_TRIG_MASK               (32'h80000000)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                                 (32'h1100)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                                 (32'h1100)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                                 (32'h1104)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                                 (32'h1104)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_R                                   (32'h1108)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_R                                   (32'h1108)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_R                                   (32'h110c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_R                                   (32'h110c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_R                                   (32'h1110)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_R                                   (32'h1110)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_R                                   (32'h1114)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_R                                   (32'h1114)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_R                                   (32'h1118)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_R                                   (32'h1118)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_R                                   (32'h111c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_R                                   (32'h111c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_R                                   (32'h1120)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_R                                   (32'h1120)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_R                                   (32'h1124)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_R                                   (32'h1124)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_R                                   (32'h1128)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_R                                   (32'h1128)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_R                                   (32'h112c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_R                                   (32'h112c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_R                                  (32'h1130)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_R                                  (32'h1130)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_R                                  (32'h1134)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_R                                  (32'h1134)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_R                                  (32'h1138)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_R                                  (32'h1138)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_R                                  (32'h113c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_R                                  (32'h113c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_R                                  (32'h1140)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_R                                  (32'h1140)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_R                                  (32'h1144)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_R                                  (32'h1144)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_R                                  (32'h1148)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_R                                  (32'h1148)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_R                                  (32'h114c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_R                                  (32'h114c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_R                                  (32'h1150)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_R                                  (32'h1150)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_R                                  (32'h1154)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_R                                  (32'h1154)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_R                                  (32'h1158)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_R                                  (32'h1158)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_R                                  (32'h115c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_R                                  (32'h115c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_R                                  (32'h1160)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_R                                  (32'h1160)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_R                                  (32'h1164)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_R                                  (32'h1164)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_R                                  (32'h1168)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_R                                  (32'h1168)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_R                                  (32'h116c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_R                                  (32'h116c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_R                                  (32'h1170)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_R                                  (32'h1170)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_R                                  (32'h1174)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_R                                  (32'h1174)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_R                                  (32'h1178)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_R                                  (32'h1178)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_R                                  (32'h117c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_R                                  (32'h117c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_R                                  (32'h1180)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_R                                  (32'h1180)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_R                                  (32'h1184)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_R                                  (32'h1184)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_R                                   (32'h1200)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_R                                   (32'h1200)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_R                                (32'h1204)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_R                                (32'h1204)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_R                               (32'h1208)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_R                               (32'h1208)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_R                               (32'h120c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_R                               (32'h120c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_R                               (32'h1210)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_R                               (32'h1210)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_R                               (32'h1214)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_R                               (32'h1214)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_R                               (32'h1218)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_R                               (32'h1218)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_R                               (32'h121c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_R                               (32'h121c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_R                               (32'h1220)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_R                               (32'h1220)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_R                               (32'h1224)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_R                               (32'h1224)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_R                               (32'h1228)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_R                               (32'h1228)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_R                               (32'h122c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_R                               (32'h122c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_R                              (32'h1230)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_R                              (32'h1230)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_R                              (32'h1234)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_R                              (32'h1234)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_R                              (32'h1238)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_R                              (32'h1238)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_R                              (32'h123c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_R                              (32'h123c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_R                              (32'h1240)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_R                              (32'h1240)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_R                              (32'h1244)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_R                              (32'h1244)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_R                              (32'h1248)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_R                              (32'h1248)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_R                              (32'h124c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_R                              (32'h124c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_R                              (32'h1250)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_R                              (32'h1250)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_R                              (32'h1254)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_R                              (32'h1254)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_R                              (32'h1258)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_R                              (32'h1258)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_R                              (32'h125c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_R                              (32'h125c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_R                              (32'h1260)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_R                              (32'h1260)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_R                              (32'h1264)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_R                              (32'h1264)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_R                              (32'h1268)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_R                              (32'h1268)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_R                              (32'h126c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_R                              (32'h126c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_R                              (32'h1270)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_R                              (32'h1270)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_R                              (32'h1274)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_R                              (32'h1274)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_R                              (32'h1278)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_R                              (32'h1278)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_R                              (32'h127c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_R                              (32'h127c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_R                              (32'h1280)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_R                              (32'h1280)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_R                              (32'h1284)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_R                              (32'h1284)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                            (32'h1300)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                            (32'h1300)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R_PULSE_LOW                  (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R_PULSE_MASK                 (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                            (32'h1304)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                            (32'h1304)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R_PULSE_LOW                  (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R_PULSE_MASK                 (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R                              (32'h1308)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R                              (32'h1308)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R                              (32'h130c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R                              (32'h130c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R                              (32'h1310)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R                              (32'h1310)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R                              (32'h1314)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R                              (32'h1314)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R                              (32'h1318)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R                              (32'h1318)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R                              (32'h131c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R                              (32'h131c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R                              (32'h1320)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R                              (32'h1320)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R                              (32'h1324)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R                              (32'h1324)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R                              (32'h1328)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R                              (32'h1328)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R                              (32'h132c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R                              (32'h132c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R                             (32'h1330)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R                             (32'h1330)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R                             (32'h1334)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R                             (32'h1334)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R                             (32'h1338)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R                             (32'h1338)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R                             (32'h133c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R                             (32'h133c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R                             (32'h1340)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R                             (32'h1340)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R                             (32'h1344)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R                             (32'h1344)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R                             (32'h1348)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R                             (32'h1348)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R                             (32'h134c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R                             (32'h134c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R                             (32'h1350)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R                             (32'h1350)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R                             (32'h1354)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R                             (32'h1354)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R                             (32'h1358)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R                             (32'h1358)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R                             (32'h135c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R                             (32'h135c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R                             (32'h1360)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R                             (32'h1360)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R                             (32'h1364)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R                             (32'h1364)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R                             (32'h1368)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R                             (32'h1368)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R                             (32'h136c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R                             (32'h136c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R                             (32'h1370)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R                             (32'h1370)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R                             (32'h1374)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R                             (32'h1374)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R                             (32'h1378)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R                             (32'h1378)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R                             (32'h137c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R                             (32'h137c)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R                             (32'h1380)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R                             (32'h1380)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R                             (32'h1384)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R                             (32'h1384)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R                              (32'h1388)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R                              (32'h1388)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_INCR_R                           (32'h138c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_INCR_R                           (32'h138c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_INCR_R_PULSE_LOW                 (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_CLPRA_MCU_RESET_REQ_INTR_COUNT_INCR_R_PULSE_MASK                (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R                          (32'h1390)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R                          (32'h1390)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R                          (32'h1394)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R                          (32'h1394)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R                          (32'h1398)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R                          (32'h1398)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R                          (32'h139c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R                          (32'h139c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R                          (32'h13a0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R                          (32'h13a0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R                          (32'h13a4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R                          (32'h13a4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R                          (32'h13a8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R                          (32'h13a8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R                          (32'h13ac)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R                          (32'h13ac)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R                          (32'h13b0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R                          (32'h13b0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R                          (32'h13b4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R                          (32'h13b4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R_PULSE_LOW                (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R_PULSE_MASK               (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R                         (32'h13b8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R                         (32'h13b8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R                         (32'h13bc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R                         (32'h13bc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R                         (32'h13c0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R                         (32'h13c0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R                         (32'h13c4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R                         (32'h13c4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R                         (32'h13c8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R                         (32'h13c8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R                         (32'h13cc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R                         (32'h13cc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R                         (32'h13d0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R                         (32'h13d0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R                         (32'h13d4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R                         (32'h13d4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R                         (32'h13d8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R                         (32'h13d8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R                         (32'h13dc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R                         (32'h13dc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R                         (32'h13e0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R                         (32'h13e0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R                         (32'h13e4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R                         (32'h13e4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R                         (32'h13e8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R                         (32'h13e8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R                         (32'h13ec)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R                         (32'h13ec)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R                         (32'h13f0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R                         (32'h13f0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R                         (32'h13f4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R                         (32'h13f4)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R                         (32'h13f8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R                         (32'h13f8)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R                         (32'h13fc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R                         (32'h13fc)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R                         (32'h1400)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R                         (32'h1400)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R                         (32'h1404)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R                         (32'h1404)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R                         (32'h1408)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R                         (32'h1408)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R                         (32'h140c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R                         (32'h140c)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R_PULSE_LOW               (0)
`define MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R_PULSE_MASK              (32'h1)


`endif