
//********************************************************************************
// SPDX-License-Identifier: Apache-2.0
// 
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//********************************************************************************

`timescale 1ps/1ps

`include "soc_address_map_defines.svh"
`include "caliptra_ss_top_tb_intc_includes.svh"

module aaxi4_interconnect(
    input logic		core_clk,	
    input logic      rst_l);

import aaxi_pkg::*;
import aaxi_pkg_xactor::*;
import aaxi_pkg_test::*;
import aaxi_pll::*;
import aaxi_pkg_caliptra_test::*;

// AXI Reset, Deassert=H, Assert=L
// bit         rst_l;
wire        ACLK;               // AXI Clock, it was generated by pll class


// low power interface
wire		   CSYSREQ;
wire		   CACTIVE;
wire		   CACTIVE_PLL;
wire		   CSYSACK;
wire		   CSYSACK_PLL;

// pll class 
// aaxi_class_pll sys_pll;

// device classes
aaxi_interconnect intc;
aaxi_device_class master[AAXI_INTC_MASTER_CNT];
aaxi_device_class slave[AAXI_INTC_SLAVE_CNT];

// device interface
// aaxi_pll_intf		ports_intf		(core_clk, rst_l, CACTIVE_PLL, CSYSREQ, CSYSACK_PLL);
aaxi_interconnect_intf	ports			(core_clk, rst_l, CACTIVE, 1'b0/*CSYSREQ*/, CSYSACK);
aaxi_intf #(.MCB_INPUT(aaxi_pkg::AAXI_MCB_INPUT),.MCB_OUTPUT(aaxi_pkg::AAXI_MCB_OUTPUT),.SCB_INPUT(aaxi_pkg::AAXI_SCB_INPUT),.SCB_OUTPUT(aaxi_pkg::AAXI_SCB_OUTPUT))mintf_arr[AAXI_INTC_MASTER_CNT-1:0]	(core_clk, rst_l, CACTIVE, 1'b0/*CSYSREQ*/, CSYSACK);
aaxi_intf #(.MCB_INPUT(aaxi_pkg::AAXI_MCB_INPUT),.MCB_OUTPUT(aaxi_pkg::AAXI_MCB_OUTPUT),.SCB_INPUT(aaxi_pkg::AAXI_SCB_INPUT),.SCB_OUTPUT(aaxi_pkg::AAXI_SCB_OUTPUT))sintf_arr[AAXI_INTC_SLAVE_CNT-1:0]	(core_clk, rst_l, CACTIVE, 1'b0/*CSYSREQ*/, CSYSACK);

/* When all CACTIVE signal of ports, mintf_arr[] and sintf_arr[] 
   are different from each other(some ports whose CACTIVE was 1,
   these ports has transaction to write or read), 
   the CACTIVE_PLL will be set 1 (can not enter low power state) */
assign CACTIVE_PLL = ((CACTIVE === 1'bx)? 1: CACTIVE);
/* When all CSYSACK signal of ports, mintf_arr[] and sintf_arr[]
   are different from each other(some ports whose CSYSACK was 1,
   these ports has transaction to write or read), 
   the CSYSACK_PLL will be set 1 (can not enter low power state) */
assign CSYSACK_PLL = ((CSYSACK === 1'bx)? 1: CSYSACK);

genvar i;
generate
    for ( i = 0; i < AAXI_INTC_MASTER_CNT; i++ ) begin : master_loop
	initial begin
	    master[i] = new($psprintf("master%0d" ,i), AAXI_MASTER, AAXI4, mintf_arr[i],, i);
	    #1;	// wait to instantiate intc bfm 
	    intc.master_ports[i].vers= master[i].vers;
	    intc.master_ports[i].ports= mintf_arr[i];
	end
    assign mintf_arr[i].CACTIVE_m = 1'b0;
    assign mintf_arr[i].CACTIVE_s = 1'b0;
    assign mintf_arr[i].CSYSACK_m = 1'b0;
    assign mintf_arr[i].CSYSACK_s = 1'b0;
    end

    for ( i = 0; i < AAXI_INTC_SLAVE_CNT; i++ ) begin: slave_loop
	initial begin
	    slave[i] = new($psprintf("slave%0d", i), AAXI_SLAVE_TO_INTERCONNECT, AAXI4, sintf_arr[i],, i);
	    #1;	// wait to instantiate intc bfm 
	    intc.slave_ports[i].vers= slave[i].vers;
	    intc.slave_ports[i].ports= sintf_arr[i];
	end
    assign sintf_arr[i].CACTIVE_m = 1'b0;
    assign sintf_arr[i].CACTIVE_s = 1'b0;
    assign sintf_arr[i].CSYSACK_m = 1'b0;
    assign sintf_arr[i].CSYSACK_s = 1'b0;
    end
endgenerate 


// bus monitor/checker0
`ifdef AVERY_ASSERT_ON

generate 
    // interfaces between Master BFMs and Interconnect slave ports
    for ( i = 0; i < AAXI_INTC_MASTER_CNT; i++ ) begin: master_mon
        aaxi_monitor_wrapper monitor(mintf_arr[i]);
        defparam monitor.VER= "AXI4";
        defparam monitor.ID_WIDTH= AAXI_ID_WIDTH;
        defparam monitor.monitor.FNAME_TRACK= {"m0"+i,"_intf.txt"};
        defparam monitor.checker0.RecMaxWaitOn= 0;
    end
    // MCU IFU, LSU, SB i/fs
    defparam master_mon[`CSS_INTC_MINTF_MCU_LSU_IDX].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    defparam master_mon[`CSS_INTC_MINTF_MCU_IFU_IDX].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    defparam master_mon[`CSS_INTC_MINTF_MCU_SB_IDX ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    // Caliptra AXI DMA, SoC BFM i/fs
    defparam master_mon[`CSS_INTC_MINTF_CPTRA_DMA_IDX].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    defparam master_mon[`CSS_INTC_MINTF_SOC_BFM_IDX  ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)

    // interfaces between Slave BFMs and Interconnect master ports
    for ( i = 0; i < AAXI_INTC_SLAVE_CNT; i++ ) begin: slave_mon
        aaxi_monitor_wrapper monitor(sintf_arr[i]);
        defparam monitor.VER= "AXI4";
        defparam monitor.ID_WIDTH= AAXI_INTC_ID_WIDTH;
        defparam monitor.monitor.FNAME_TRACK= {"s0"+i,"_intf.txt"};
        defparam monitor.checker0.RecMaxWaitOn= 0;
    end
    // NC, MCU ROM, FC PRIM (NC)
    defparam slave_mon[`CSS_INTC_SINTF_NC0_IDX    ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    defparam slave_mon[`CSS_INTC_SINTF_MCU_ROM_IDX].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    defparam slave_mon[`CSS_INTC_SINTF_NC1_IDX    ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH; // set DATA BUS WIDTH to match interconnect native width
    // I3C, Caliptra SoC IFC, MCI, FC, LCC
    defparam slave_mon[`CSS_INTC_SINTF_I3C_IDX          ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    defparam slave_mon[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    defparam slave_mon[`CSS_INTC_SINTF_MCI_IDX          ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    defparam slave_mon[`CSS_INTC_SINTF_FC_IDX           ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    defparam slave_mon[`CSS_INTC_SINTF_LCC_IDX          ].monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH/2; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        
endgenerate 

// instantiates monitor/protocol checker0 for default slave interface
assign ports.default_slave_intf.CACTIVE_m = 1'b0;
assign ports.default_slave_intf.CACTIVE_s = 1'b0;
assign ports.default_slave_intf.CSYSACK_m = 1'b0;
assign ports.default_slave_intf.CSYSACK_s = 1'b0;
aaxi_monitor_wrapper def_monitor(ports.default_slave_intf);
defparam def_monitor.VER= "AXI4";
defparam def_monitor.ID_WIDTH= AAXI_INTC_ID_WIDTH;
defparam def_monitor.BUS_DATA_WIDTH= AAXI_DATA_WIDTH;    // set DATA BUS WIDTH
defparam def_monitor.checker0.RecMaxWaitOn= 0;
defparam def_monitor.monitor.FNAME_TRACK= "default_slave_intf.txt";

`endif

// instance device classes

int j, depth2;
aaxi_priority_tier_type priority_master;


initial begin
    #0;
    intc = new("intc", AAXI_INTERCONNECT,, ports);
    // PLL class, instantiates clock generator
    // sys_pll = new("Avery_pll", ports_intf);
    #0;

    for (int i = 0; i < AAXI_INTC_MASTER_CNT; i++) begin
        // instantiates Master BFMs
        master[i].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        master[i].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        master[i].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        master[i].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        master[i].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        master[i].cfg_info.passive_mode= 1;       //-- changed to put master to passive mode
        // master[i].cfg_info.id_width=3;
`ifdef FOUR_OUTSTANDING
        master[i].cfg_info.total_outstanding_depth = 4;
        master[i].cfg_info.id_outstanding_depth = 4;
`else
        master[i].cfg_info.total_outstanding_depth = 1;
        master[i].cfg_info.id_outstanding_depth = 1;
`endif
        master[i].cfg_info.no_overlap_allow = 0;
`ifdef UNALIGNED_WSTRB_ONLY
        master[i].cfg_info.unaligned_transfer_addr = 1;
`endif
`ifdef DEFAULT_HIGH
        master[i].cfg_info.bready_default = 1;
        master[i].cfg_info.rready_default = 1;
`endif
    end

    master[`CSS_INTC_MINTF_MCU_LSU_IDX].  cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width
    master[`CSS_INTC_MINTF_MCU_IFU_IDX].  cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width
    master[`CSS_INTC_MINTF_MCU_SB_IDX].   cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width
    master[`CSS_INTC_MINTF_CPTRA_DMA_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
    master[`CSS_INTC_MINTF_SOC_BFM_IDX].  cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)

    wait (slave[0] != null);
    for (int i=0; i<AAXI_INTC_SLAVE_CNT; i++) begin
        // instantiates Slave BFMs
        slave[i].cfg_info.passive_mode= 1; 
        slave[i].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[i].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[i].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[i].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[i].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        // slave[i].add_fifo(64'habcc+i*64'h100_0000, 4);
        // slave[i].add_fifo(64'ha000_0000+i*64'h100_0000, 4);
        // slave[i].add_fifo(64'hb000_0001+i*64'h100_0000, 4);
        // slave[i].cfg_info.fifo_address[0] = 64'hc000_0000;
        // slave[i].cfg_info.fifo_limit[0] = 64'hc000_1000;
`ifdef FOUR_OUTSTANDING
        slave[i].cfg_info.total_outstanding_depth = 4;
        slave[i].cfg_info.id_outstanding_depth = 4;
`else
        slave[i].cfg_info.total_outstanding_depth = 1;
        slave[i].cfg_info.id_outstanding_depth = 1;
`endif
`ifdef DEFAULT_HIGH
        slave[i].cfg_info.awready_default = 1;
        slave[i].cfg_info.dwready_default = 1;
        slave[i].cfg_info.arready_default = 1;
`endif
    end
        //-- Not Connected
        slave[`CSS_INTC_SINTF_NC0_IDX].cfg_info.base_address[0]  = 64'h1000_0000;
        slave[`CSS_INTC_SINTF_NC0_IDX].cfg_info.limit_address[0] = 64'h1000_FFFF;
        slave[`CSS_INTC_SINTF_NC0_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width

        //-- I3C
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.passive_mode = 1;
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.base_address[0] = 64'h2000_4000;
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.limit_address[0] = 64'h2000_4FFF;
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_I3C_IDX].cfg_info.id_outstanding_depth = 4;

        //-- MCU ROM MACRO / MCI_TOP 2nd instance
        slave[`CSS_INTC_SINTF_MCU_ROM_IDX].cfg_info.base_address[0] = {32'h0, 32'h8000_0000};
        slave[`CSS_INTC_SINTF_MCU_ROM_IDX].cfg_info.limit_address[0] = {32'h0, 32'h80FF_FFFF};
        slave[`CSS_INTC_SINTF_MCU_ROM_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width

        //-- Caliptra SoC IFC Sub
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.passive_mode= 1; 
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.base_address[0] = 64'(`SOC_MBOX_CSR_BASE_ADDR);
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.limit_address[0] = 64'(`SOC_MBOX_CSR_BASE_ADDR) + 64'h2_0000; // FIXME hardcoded to match the soc_ifc limit
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.default_fifo_depth = 4096; // Reasonable cap at max AXI burst lengh of 4KiB
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.fifo_address[0] = 64'(`SOC_MBOX_CSR_MBOX_DATAIN);
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.fifo_limit[0] = 64'(`SOC_MBOX_CSR_MBOX_DATAOUT);
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.fifo_address[1] = 64'(`SOC_SHA512_ACC_CSR_DATAIN);
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.fifo_limit[1] = 64'(`SOC_SHA512_ACC_CSR_DATAIN);
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_CPTRA_SOC_IFC_IDX].cfg_info.id_outstanding_depth = 4;

        //-- MCI
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.passive_mode= 1; 
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.base_address[0]  = {32'h0, `SOC_MCI_TOP_MCI_REG_BASE_ADDR}; //64'h2100_0000;
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.limit_address[0] = {32'h0, `SOC_MCI_TOP_MCU_SRAM_END_ADDR}; // Always the last address in MCU
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_MCI_IDX].cfg_info.id_outstanding_depth = 4;

        //-- Fuse Controller Core AXI 
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.passive_mode = 1; 
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.base_address[0] = {32'h0, `SOC_OTP_CTRL_BASE_ADDR}; //64'h7000_0000;
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.limit_address[0] = {32'h0, `SOC_OTP_CTRL_BASE_ADDR} + 'h1FF; //64'h7000_01FF;
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_FC_IDX].cfg_info.id_outstanding_depth = 4;

        //-- Fuse Controller Prim AXI (not connected)
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.passive_mode = 1; 
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.base_address[0] = 64'h7000_0200;
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.limit_address[0] = 64'h7000_03FF;
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 3; // set DATA BUS WIDTH to match interconnect native width
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_NC1_IDX].cfg_info.id_outstanding_depth = 4;

        //-- Life-cycle Controller Core AXI 
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.passive_mode = 1; 
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.opt_awuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.opt_aruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.opt_ruser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.opt_wuser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.opt_buser_enable = 1; // optional, axi4_interconn_routings.sv need it
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.base_address[0] = {32'h0, `SOC_LC_CTRL_BASE_ADDR}; //64'h7000_0400;
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.limit_address[0] = {32'h0, `SOC_LC_CTRL_BASE_ADDR} + 'h5FF;// 64'h7000_05FF;
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.data_bus_bytes = AAXI_DATA_WIDTH >> 4; // set DATA BUS WIDTH to interconnect native width / 2 (32b)
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.total_outstanding_depth = 4;
        slave[`CSS_INTC_SINTF_LCC_IDX].cfg_info.id_outstanding_depth = 4;



//#1;
//do not sure what feature of #1
    // connect devices to the Interconnect
    for (int i=0; i<AAXI_INTC_MASTER_CNT; i++) begin
	j = (i+2)%3;
	priority_master = aaxi_priority_tier_type'(j);
	master[i].cfg_info.ms_priority= priority_master;
	master[i].cfg_info.copy_partial_fields(intc.master_ports[i].cfg_info);
    end
    for (int i=0; i<AAXI_INTC_SLAVE_CNT; i++) begin
	slave[i].cfg_info.copy_partial_fields(intc.slave_ports[i].cfg_info);
    end

    depth2= 1;
`ifdef INTERCONNECT_PORT_INTERLEAVE_FOUR
    depth2= 4;
`endif
    for (int i=0; i < AAXI_INTC_MASTER_CNT; i++) begin
`ifdef INTERCONNECT_DEFAULT_LOW
	// set the default ready of intc ports as zero
	intc.set_port_default_ready(i, 1, AAXI_ALL_READY, 0);
`endif

	// set the write/read interleave depth of Interconnect slave/master ports as four
	intc.set_port_interleave_depth(i, 1, depth2);

`ifdef INTERCONNECT_BUS_BUFFER_SIZE_FOUR
	// set the buffer size of data/resp buses inside Interconnect
	intc.set_port_bus_buffer_size(AAXI_BUS_TYPE_READ_DATA, 4, i);
	intc.set_port_bus_buffer_size(AAXI_BUS_TYPE_WRITE_RESP, 4, i);
`endif
	end


    for (int i=0; i < AAXI_INTC_SLAVE_CNT; i++) begin
`ifdef INTERCONNECT_DEFAULT_LOW
	// set the default ready of intc ports as zero
	intc.set_port_default_ready(i, 0, AAXI_ALL_READY, 0);
`endif

	// set the write/read interleave depth of Interconnect slave/master ports as four
	intc.set_port_interleave_depth(i, 0, depth2);

`ifdef INTERCONNECT_BUS_BUFFER_SIZE_FOUR
	// set the buffer size of data buses inside Interconnect
	intc.set_port_bus_buffer_size(AAXI_BUS_TYPE_WRITE_DATA, 4, i);
`endif
	end

`ifdef INTERCONNECT_BUS_BUFFER_SIZE_FOUR
    // set the buffer size of write/read address bus inside Interconnect
    intc.set_port_bus_buffer_size(AAXI_BUS_TYPE_WRITE_ADDR, 4);
    intc.set_port_bus_buffer_size(AAXI_BUS_TYPE_READ_ADDR, 4);
`endif
    end

    //task automatic start_test(aaxi_test_base test);
    task automatic start_test(aaxi_test_caliptra_ss test);
        aaxi_pkg_test::aaxi_test_select(test.test_name);
        test.master0= master[0];
        test.master1= master[1];
        test.master2= master[2];
        test.master3= master[3];
        for (int i=0; i< AAXI_INTC_MASTER_CNT; i++) begin
        test.ms_bfms.push_back(master[i]);
    `ifdef PASSIVE_MASTER
        test.psv_ms_bfms.push_back(passive_master[i]);
    `endif
        end

        // initial memory value to be 0 for data comparision on Slave BFM 
        slave[0].set("mem_uninitialized_value", 0);
        slave[1].set("mem_uninitialized_value", 0);
        slave[2].set("mem_uninitialized_value", 0);
        slave[3].set("mem_uninitialized_value", 0);
        slave[4].set("mem_uninitialized_value", 0);
        slave[5].set("mem_uninitialized_value", 0);
        slave[6].set("mem_uninitialized_value", 0);
        slave[7].set("mem_uninitialized_value", 0);


        test.slave0= slave[0];
        test.slave1= slave[1];
        test.slave2= slave[2];
        test.slave3= slave[3];
        test.slave4= slave[4];
        test.slave5= slave[5];
        test.slave6= slave[6];
        test.slave7= slave[7];

        for (int i=0; i< AAXI_INTC_SLAVE_CNT; i++)
            test.slv_bfms.push_back(slave[i]);

        test.itc_bfm= intc;
    `ifdef PASSIVE_ITC
        test.psv_itc_bfm= passive_intc;
    `endif
        test.run();
    endtask
endmodule

