// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//



`include "mci_common_tasks.svh"
`include "mci_mcu_trace_buffer_mon.svh"
`include "smoke_test_mcu_sram_execution_region.svh"
`include "smoke_test_mcu_sram_debug_stress.svh"
`include "smoke_test_mcu_trace_buffer.svh"
`include "mcu_mbox_soc_agent_write_fw_image.svh"
`include "smoke_test_mcu_trace_buffer_no_debug.svh"
`include "smoke_test_mci_soc_config_disable.svh"
`include "smoke_test_mci_soc_config_always_enable.svh"
`include "smoke_test_mci_soc_config_diff_mcu.svh"
