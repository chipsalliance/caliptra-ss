
`ifndef CPTRA_SS_INCLUDES_SVH
`define CPTRA_SS_INCLUDES_SVH


parameter CPTRA_SS_MCU_USER_WIDTH = 32;

parameter CALIPTRA_CORE_AXI_USER_ID =          32'h0;
parameter MCU_AXI_USER_ID           =          32'h1;

`endif // CPTRA_SS_INCLUDES_SVH