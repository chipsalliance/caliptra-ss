//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in register_test.
// It uses the UVM built in register test.  Specific UVM built-in tests can be
// selected in the body task.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

class register_test_sequence extends fuse_ctrl_bench_sequence_base;

  `uvm_object_utils( register_test_sequence );


  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end

  function new(string name = "" );
    super.new(name);
  endfunction

  // ****************************************************************************
  virtual task body();

    // Reset the DUT
    fork
      // pragma uvmf custom register_test_reset begin
      // UVMF_CHANGE_ME 
      // Select the desired wait_for_reset or provide custom mechanism.
      // fork-join for this code block may be unnecessary based on your situation.
      fuse_ctrl_rst_in_agent_config.wait_for_reset();
      fuse_ctrl_rst_out_agent_config.wait_for_reset();
      fuse_ctrl_core_axi_write_in_if_agent_config.wait_for_reset();
      fuse_ctrl_core_axi_write_out_if_agent_config.wait_for_reset();
      fuse_ctrl_prim_axi_write_in_if_agent_config.wait_for_reset();
      fuse_ctrl_prim_axi_write_out_if_agent_config.wait_for_reset();
      fuse_ctrl_core_axi_read_in_if_agent_config.wait_for_reset();
      fuse_ctrl_core_axi_read_out_if_agent_config.wait_for_reset();
      fuse_ctrl_prim_axi_read_in_if_agent_config.wait_for_reset();
      fuse_ctrl_prim_axi_read_out_if_agent_config.wait_for_reset();
      fuse_ctrl_secreg_axi_read_in_if_agent_config.wait_for_reset();
      fuse_ctrl_secreg_axi_read_out_if_agent_config.wait_for_reset();
      fuse_ctrl_lc_otp_in_if_agent_config.wait_for_reset();
      fuse_ctrl_lc_otp_out_if_agent_config.wait_for_reset();
      fuse_ctrl_in_if_agent_config.wait_for_reset();
      fuse_ctrl_out_if_agent_config.wait_for_reset();
      // pragma uvmf custom register_test_reset end
    join

      // pragma uvmf custom register_test_setup begin
      // UVMF_CHANGE_ME perform potentially necessary operations before running the sequence.
      // pragma uvmf custom register_test_setup end

    // pragma uvmf custom register_test_operation begin
    // UVMF_CHANGE_ME Perform your custom register test
    // pragma uvmf custom register_test_operation end

  endtask

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

