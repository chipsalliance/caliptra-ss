
`ifndef CPTRA_SS_INCLUDES_SVH
`define CPTRA_SS_INCLUDES_SVH


parameter CPTRA_SS_MCU_USER_WIDTH = 32;

`endif // CPTRA_SS_INCLUDES_SVH