`include "config_defines_mcu.svh"
