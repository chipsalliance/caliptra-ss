// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

`include "cptra_ss_i3c_core_defines.svh"
`include "cptra_ss_i3c_core_base_test.svh"
`include "i3c_reg_rd_wr.svh"
`include "i3c_sboot.svh"
`include "ai3ct_ext_basic.svh"
