`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 03/21/2023 11:49:47 AM
// Design Name:
// Module Name: caliptra_package_top
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments: Vivado does not support using a SystemVerilog as the top level file in an package.
//
//////////////////////////////////////////////////////////////////////////////////

`default_nettype wire

`define CALIPTRA_APB_ADDR_WIDTH      32 // bit-width APB address
`define CALIPTRA_APB_DATA_WIDTH      32 // bit-width APB data

module caliptra_package_axi_top (
    input wire core_clk,
    input wire i3c_clk,

    input wire axi_i3c_scl_t,
    input wire axi_i3c_scl_o,
    input wire axi_i3c_scl_pullup_en,
    input wire axi_i3c_sda_t,
    input wire axi_i3c_sda_o,
    input wire axi_i3c_sda_pullup_en,
    // I3C signals back to AXI I3C
    output wire SCL,
    output wire SDA,

    // Caliptra AXI Interface
    input  wire [31:0] S_AXI_CALIPTRA_AWADDR,
    input  wire [1:0] S_AXI_CALIPTRA_AWBURST,
    input  wire [2:0] S_AXI_CALIPTRA_AWSIZE,
    input  wire [7:0] S_AXI_CALIPTRA_AWLEN,
    input  wire [31:0] S_AXI_CALIPTRA_AWUSER,
    input  wire [15:0] S_AXI_CALIPTRA_AWID,
    input  wire S_AXI_CALIPTRA_AWLOCK,
    input  wire S_AXI_CALIPTRA_AWVALID,
    output wire S_AXI_CALIPTRA_AWREADY,
    // W
    input  wire [31:0] S_AXI_CALIPTRA_WDATA,
    input  wire [3:0] S_AXI_CALIPTRA_WSTRB,
    input  wire S_AXI_CALIPTRA_WVALID,
    output wire S_AXI_CALIPTRA_WREADY,
    input  wire S_AXI_CALIPTRA_WLAST,
    // B
    output wire [1:0] S_AXI_CALIPTRA_BRESP,
    output wire [15:0] S_AXI_CALIPTRA_BID,
    output wire S_AXI_CALIPTRA_BVALID,
    input  wire S_AXI_CALIPTRA_BREADY,
    // AR
    input  wire [31:0] S_AXI_CALIPTRA_ARADDR,
    input  wire [1:0] S_AXI_CALIPTRA_ARBURST,
    input  wire [2:0] S_AXI_CALIPTRA_ARSIZE,
    input  wire [7:0] S_AXI_CALIPTRA_ARLEN,
    input  wire [31:0] S_AXI_CALIPTRA_ARUSER,
    input  wire [15:0] S_AXI_CALIPTRA_ARID,
    input  wire S_AXI_CALIPTRA_ARLOCK,
    input  wire S_AXI_CALIPTRA_ARVALID,
    output wire S_AXI_CALIPTRA_ARREADY,
    // R
    output wire [31:0] S_AXI_CALIPTRA_RDATA,
    output wire [1:0] S_AXI_CALIPTRA_RRESP,
    output wire [15:0] S_AXI_CALIPTRA_RID,
    output wire S_AXI_CALIPTRA_RLAST,
    output wire S_AXI_CALIPTRA_RVALID,
    input  wire S_AXI_CALIPTRA_RREADY,

    // Caliptra M_AXI Interface
    output  wire [31:0] M_AXI_CALIPTRA_AWADDR,
    output  wire [1:0] M_AXI_CALIPTRA_AWBURST,
    output  wire [2:0] M_AXI_CALIPTRA_AWSIZE,
    output  wire [7:0] M_AXI_CALIPTRA_AWLEN,
    output  wire [31:0] M_AXI_CALIPTRA_AWUSER,
    output  wire [15:0] M_AXI_CALIPTRA_AWID,
    output  wire M_AXI_CALIPTRA_AWLOCK,
    output  wire M_AXI_CALIPTRA_AWVALID,
    input wire M_AXI_CALIPTRA_AWREADY,
    // W
    output  wire [31:0] M_AXI_CALIPTRA_WDATA,
    output  wire [3:0] M_AXI_CALIPTRA_WSTRB,
    output  wire M_AXI_CALIPTRA_WVALID,
    input wire M_AXI_CALIPTRA_WREADY,
    output  wire M_AXI_CALIPTRA_WLAST,
    // B
    input wire [1:0] M_AXI_CALIPTRA_BRESP,
    input wire  [15:0] M_AXI_CALIPTRA_BID,
    input wire M_AXI_CALIPTRA_BVALID,
    output  wire M_AXI_CALIPTRA_BREADY,
    // AR
    output  wire [31:0] M_AXI_CALIPTRA_ARADDR,
    output  wire [1:0] M_AXI_CALIPTRA_ARBURST,
    output  wire [2:0] M_AXI_CALIPTRA_ARSIZE,
    output  wire [7:0] M_AXI_CALIPTRA_ARLEN,
    output  wire [31:0] M_AXI_CALIPTRA_ARUSER,
    output  wire [15:0] M_AXI_CALIPTRA_ARID,
    output  wire M_AXI_CALIPTRA_ARLOCK,
    output  wire M_AXI_CALIPTRA_ARVALID,
    input wire M_AXI_CALIPTRA_ARREADY,
    // R
    input wire [31:0] M_AXI_CALIPTRA_RDATA,
    input wire [1:0] M_AXI_CALIPTRA_RRESP,
    input wire [15:0] M_AXI_CALIPTRA_RID,
    input wire M_AXI_CALIPTRA_RLAST,
    input wire M_AXI_CALIPTRA_RVALID,
    output  wire M_AXI_CALIPTRA_RREADY,

    // MCI S_AXI Interface
    input  wire [31:0] S_AXI_MCI_AWADDR,
    input  wire [1:0] S_AXI_MCI_AWBURST,
    input  wire [2:0] S_AXI_MCI_AWSIZE,
    input  wire [7:0] S_AXI_MCI_AWLEN,
    input  wire [31:0] S_AXI_MCI_AWUSER,
    input  wire [15:0] S_AXI_MCI_AWID,
    input  wire S_AXI_MCI_AWLOCK,
    input  wire S_AXI_MCI_AWVALID,
    output wire S_AXI_MCI_AWREADY,
    // W
    input  wire [31:0] S_AXI_MCI_WDATA,
    input  wire [3:0] S_AXI_MCI_WSTRB,
    input  wire S_AXI_MCI_WVALID,
    output wire S_AXI_MCI_WREADY,
    input  wire S_AXI_MCI_WLAST,
    // B
    output wire [1:0] S_AXI_MCI_BRESP,
    output wire [15:0] S_AXI_MCI_BID,
    output wire S_AXI_MCI_BVALID,
    input  wire S_AXI_MCI_BREADY,
    // AR
    input  wire [31:0] S_AXI_MCI_ARADDR,
    input  wire [1:0] S_AXI_MCI_ARBURST,
    input  wire [2:0] S_AXI_MCI_ARSIZE,
    input  wire [7:0] S_AXI_MCI_ARLEN,
    input  wire [31:0] S_AXI_MCI_ARUSER,
    input  wire [15:0] S_AXI_MCI_ARID,
    input  wire S_AXI_MCI_ARLOCK,
    input  wire S_AXI_MCI_ARVALID,
    output wire S_AXI_MCI_ARREADY,
    // R
    output wire [31:0] S_AXI_MCI_RDATA,
    output wire [1:0] S_AXI_MCI_RRESP,
    output wire [15:0] S_AXI_MCI_RID,
    output wire S_AXI_MCI_RLAST,
    output wire S_AXI_MCI_RVALID,
    input  wire S_AXI_MCI_RREADY,

    // MCI ROM S_AXI Interface
    input  wire [31:0] S_AXI_MCU_ROM_AWADDR,
    input  wire [1:0] S_AXI_MCU_ROM_AWBURST,
    input  wire [2:0] S_AXI_MCU_ROM_AWSIZE,
    input  wire [7:0] S_AXI_MCU_ROM_AWLEN,
    input  wire [31:0] S_AXI_MCU_ROM_AWUSER,
    input  wire [15:0] S_AXI_MCU_ROM_AWID,
    input  wire S_AXI_MCU_ROM_AWLOCK,
    input  wire S_AXI_MCU_ROM_AWVALID,
    output wire S_AXI_MCU_ROM_AWREADY,
    // W
    input  wire [63:0] S_AXI_MCU_ROM_WDATA,
    input  wire [7:0] S_AXI_MCU_ROM_WSTRB,
    input  wire S_AXI_MCU_ROM_WVALID,
    output wire S_AXI_MCU_ROM_WREADY,
    input  wire S_AXI_MCU_ROM_WLAST,
    // B
    output wire [1:0] S_AXI_MCU_ROM_BRESP,
    output wire [15:0] S_AXI_MCU_ROM_BID,
    output wire S_AXI_MCU_ROM_BVALID,
    input  wire S_AXI_MCU_ROM_BREADY,
    // AR
    input  wire [31:0] S_AXI_MCU_ROM_ARADDR,
    input  wire [1:0] S_AXI_MCU_ROM_ARBURST,
    input  wire [2:0] S_AXI_MCU_ROM_ARSIZE,
    input  wire [7:0] S_AXI_MCU_ROM_ARLEN,
    input  wire [31:0] S_AXI_MCU_ROM_ARUSER,
    input  wire [15:0] S_AXI_MCU_ROM_ARID,
    input  wire S_AXI_MCU_ROM_ARLOCK,
    input  wire S_AXI_MCU_ROM_ARVALID,
    output wire S_AXI_MCU_ROM_ARREADY,
    // R
    output wire [63:0] S_AXI_MCU_ROM_RDATA,
    output wire [1:0] S_AXI_MCU_ROM_RRESP,
    output wire [15:0] S_AXI_MCU_ROM_RID,
    output wire S_AXI_MCU_ROM_RLAST,
    output wire S_AXI_MCU_ROM_RVALID,
    input  wire S_AXI_MCU_ROM_RREADY,

    // MCI M_AXI Interface
    output  wire [31:0] M_AXI_MCI_AWADDR,
    output  wire [1:0] M_AXI_MCI_AWBURST,
    output  wire [2:0] M_AXI_MCI_AWSIZE,
    output  wire [7:0] M_AXI_MCI_AWLEN,
    output  wire [31:0] M_AXI_MCI_AWUSER,
    output  wire [15:0] M_AXI_MCI_AWID,
    output  wire M_AXI_MCI_AWLOCK,
    output  wire M_AXI_MCI_AWVALID,
    input wire M_AXI_MCI_AWREADY,
    // W
    output  wire [31:0] M_AXI_MCI_WDATA,
    output  wire [3:0] M_AXI_MCI_WSTRB,
    output  wire M_AXI_MCI_WVALID,
    input wire M_AXI_MCI_WREADY,
    output  wire M_AXI_MCI_WLAST,
    // B
    input wire [1:0] M_AXI_MCI_BRESP,
    input wire [15:0] M_AXI_MCI_BID,
    input wire M_AXI_MCI_BVALID,
    output  wire M_AXI_MCI_BREADY,
    // AR
    output  wire [31:0] M_AXI_MCI_ARADDR,
    output  wire [1:0] M_AXI_MCI_ARBURST,
    output  wire [2:0] M_AXI_MCI_ARSIZE,
    output  wire [7:0] M_AXI_MCI_ARLEN,
    output  wire [31:0] M_AXI_MCI_ARUSER,
    output  wire [15:0] M_AXI_MCI_ARID,
    output  wire M_AXI_MCI_ARLOCK,
    output  wire M_AXI_MCI_ARVALID,
    input wire M_AXI_MCI_ARREADY,
    // R
    input wire [31:0] M_AXI_MCI_RDATA,
    input wire [1:0] M_AXI_MCI_RRESP,
    input wire [15:0] M_AXI_MCI_RID,
    input wire M_AXI_MCI_RLAST,
    input wire M_AXI_MCI_RVALID,
    output  wire M_AXI_MCI_RREADY,


    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_LSU_AWVALID,
    input  wire                      M_AXI_MCU_LSU_AWREADY,
    output wire [18:0]              M_AXI_MCU_LSU_AWID,
    output wire [              31:0] M_AXI_MCU_LSU_AWADDR,
    output wire [               3:0] M_AXI_MCU_LSU_AWREGION,
    output wire [               7:0] M_AXI_MCU_LSU_AWLEN,
    output wire [               2:0] M_AXI_MCU_LSU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_AWBURST,
    output wire                      M_AXI_MCU_LSU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_AWPROT,
    output wire [               3:0] M_AXI_MCU_LSU_AWQOS,

    output wire                      M_AXI_MCU_LSU_WVALID,
    input  wire                      M_AXI_MCU_LSU_WREADY,
    output wire [63:0]               M_AXI_MCU_LSU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_LSU_WSTRB,
    output wire                      M_AXI_MCU_LSU_WLAST,

    input  wire                      M_AXI_MCU_LSU_BVALID,
    output wire                      M_AXI_MCU_LSU_BREADY,
    input  wire [               1:0] M_AXI_MCU_LSU_BRESP,
    input  wire [18:0]              M_AXI_MCU_LSU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_LSU_ARVALID,
    input  wire                      M_AXI_MCU_LSU_ARREADY,
    output wire [18:0]              M_AXI_MCU_LSU_ARID,
    output wire [              31:0] M_AXI_MCU_LSU_ARADDR,
    output wire [               3:0] M_AXI_MCU_LSU_ARREGION,
    output wire [               7:0] M_AXI_MCU_LSU_ARLEN,
    output wire [               2:0] M_AXI_MCU_LSU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_ARBURST,
    output wire                      M_AXI_MCU_LSU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_ARPROT,
    output wire [               3:0] M_AXI_MCU_LSU_ARQOS,

    input  wire                      M_AXI_MCU_LSU_RVALID,
    output wire                      M_AXI_MCU_LSU_RREADY,
    input  wire [18:0]              M_AXI_MCU_LSU_RID,
    input  wire [              63:0] M_AXI_MCU_LSU_RDATA,
    input  wire [               1:0] M_AXI_MCU_LSU_RRESP,
    input  wire                      M_AXI_MCU_LSU_RLAST,

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_IFU_AWVALID,
    input  wire                      M_AXI_MCU_IFU_AWREADY,
    output wire [18:0]              M_AXI_MCU_IFU_AWID,
    output wire [              31:0] M_AXI_MCU_IFU_AWADDR,
    output wire [               3:0] M_AXI_MCU_IFU_AWREGION,
    output wire [               7:0] M_AXI_MCU_IFU_AWLEN,
    output wire [               2:0] M_AXI_MCU_IFU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_AWBURST,
    output wire                      M_AXI_MCU_IFU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_AWPROT,
    output wire [               3:0] M_AXI_MCU_IFU_AWQOS,

    output wire                      M_AXI_MCU_IFU_WVALID,
    input  wire                      M_AXI_MCU_IFU_WREADY,
    output wire [63:0]               M_AXI_MCU_IFU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_IFU_WSTRB,
    output wire                      M_AXI_MCU_IFU_WLAST,

    input  wire                      M_AXI_MCU_IFU_BVALID,
    output wire                      M_AXI_MCU_IFU_BREADY,
    input  wire [               1:0] M_AXI_MCU_IFU_BRESP,
    input  wire [18:0]              M_AXI_MCU_IFU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_IFU_ARVALID,
    input  wire                      M_AXI_MCU_IFU_ARREADY,
    output wire [18:0]              M_AXI_MCU_IFU_ARID,
    output wire [              31:0] M_AXI_MCU_IFU_ARADDR,
    output wire [               3:0] M_AXI_MCU_IFU_ARREGION,
    output wire [               7:0] M_AXI_MCU_IFU_ARLEN,
    output wire [               2:0] M_AXI_MCU_IFU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_ARBURST,
    output wire                      M_AXI_MCU_IFU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_ARPROT,
    output wire [               3:0] M_AXI_MCU_IFU_ARQOS,

    input  wire                      M_AXI_MCU_IFU_RVALID,
    output wire                      M_AXI_MCU_IFU_RREADY,
    input  wire [18:0]              M_AXI_MCU_IFU_RID,
    input  wire [              63:0] M_AXI_MCU_IFU_RDATA,
    input  wire [               1:0] M_AXI_MCU_IFU_RRESP,
    input  wire                      M_AXI_MCU_IFU_RLAST,

    //-------------------------- SB AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_SB_AWVALID,
    input  wire                      M_AXI_MCU_SB_AWREADY,
    output wire [18:0]               M_AXI_MCU_SB_AWID,
    output wire [              31:0] M_AXI_MCU_SB_AWADDR,
    output wire [               3:0] M_AXI_MCU_SB_AWREGION,
    output wire [               7:0] M_AXI_MCU_SB_AWLEN,
    output wire [               2:0] M_AXI_MCU_SB_AWSIZE,
    output wire [               1:0] M_AXI_MCU_SB_AWBURST,
    output wire                      M_AXI_MCU_SB_AWLOCK,
    output wire [               3:0] M_AXI_MCU_SB_AWCACHE,
    output wire [               2:0] M_AXI_MCU_SB_AWPROT,
    output wire [               3:0] M_AXI_MCU_SB_AWQOS,

    output wire                      M_AXI_MCU_SB_WVALID,
    input  wire                      M_AXI_MCU_SB_WREADY,
    output wire [63:0]               M_AXI_MCU_SB_WDATA,
    output wire [ 7:0]               M_AXI_MCU_SB_WSTRB,
    output wire                      M_AXI_MCU_SB_WLAST,

    input  wire                      M_AXI_MCU_SB_BVALID,
    output wire                      M_AXI_MCU_SB_BREADY,
    input  wire [               1:0] M_AXI_MCU_SB_BRESP,
    input  wire [18:0]               M_AXI_MCU_SB_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_SB_ARVALID,
    input  wire                      M_AXI_MCU_SB_ARREADY,
    output wire [18:0]               M_AXI_MCU_SB_ARID,
    output wire [              31:0] M_AXI_MCU_SB_ARADDR,
    output wire [               3:0] M_AXI_MCU_SB_ARREGION,
    output wire [               7:0] M_AXI_MCU_SB_ARLEN,
    output wire [               2:0] M_AXI_MCU_SB_ARSIZE,
    output wire [               1:0] M_AXI_MCU_SB_ARBURST,
    output wire                      M_AXI_MCU_SB_ARLOCK,
    output wire [               3:0] M_AXI_MCU_SB_ARCACHE,
    output wire [               2:0] M_AXI_MCU_SB_ARPROT,
    output wire [               3:0] M_AXI_MCU_SB_ARQOS,

    input  wire                      M_AXI_MCU_SB_RVALID,
    output wire                      M_AXI_MCU_SB_RREADY,
    input  wire [18:0]               M_AXI_MCU_SB_RID,
    input  wire [              63:0] M_AXI_MCU_SB_RDATA,
    input  wire [               1:0] M_AXI_MCU_SB_RRESP,
    input  wire                      M_AXI_MCU_SB_RLAST,

    // I3C
    input	wire                      S_AXI_I3C_AWVALID,
    output	wire                      S_AXI_I3C_AWREADY,
    input	wire [31:0]               S_AXI_I3C_AWADDR,
    input	wire [2:0]                S_AXI_I3C_AWPROT,
    input	wire                      S_AXI_I3C_WVALID,
    output	wire                      S_AXI_I3C_WREADY,
    input	wire [31:0]               S_AXI_I3C_WDATA,
    input	wire [3:0]                S_AXI_I3C_WSTRB,
    output	wire                      S_AXI_I3C_BVALID,
    input	wire                      S_AXI_I3C_BREADY,
    output	wire [1:0]                S_AXI_I3C_BRESP,
    input	wire                      S_AXI_I3C_ARVALID,
    output	wire                      S_AXI_I3C_ARREADY,
    input	wire [31:0]               S_AXI_I3C_ARADDR,
    input	wire [2:0]                S_AXI_I3C_ARPROT,
    output	wire                      S_AXI_I3C_RVALID,
    input	wire                      S_AXI_I3C_RREADY,
    output	wire [31:0]               S_AXI_I3C_RDATA,
    output	wire [1:0]                S_AXI_I3C_RRESP,
    
    input wire [1:0] S_AXI_I3C_ARBURST,
    input wire [2:0] S_AXI_I3C_ARSIZE,
    input wire [7:0] S_AXI_I3C_ARLEN,
    input wire [31:0] S_AXI_I3C_ARUSER,
    input wire [18:0] S_AXI_I3C_ARID,
    input wire S_AXI_I3C_ARLOCK,
    output wire [18:0]           S_AXI_I3C_RID,
    output wire                   S_AXI_I3C_RLAST,
    input wire [             1:0] S_AXI_I3C_AWBURST,
    input wire [             2:0] S_AXI_I3C_AWSIZE,
    input wire [             7:0] S_AXI_I3C_AWLEN,
    input wire [31:0] S_AXI_I3C_AWUSER,
    input wire [18:0] S_AXI_I3C_AWID,
    input wire                    S_AXI_I3C_AWLOCK,
    input  wire                  S_AXI_I3C_WLAST,
    output wire [18:0] S_AXI_I3C_BID,

    // LCC
    input	wire                      S_AXI_LCC_AWVALID,
    output	wire                      S_AXI_LCC_AWREADY,
    input	wire [31:0]               S_AXI_LCC_AWADDR,
    input	wire [2:0]                S_AXI_LCC_AWPROT,
    input	wire                      S_AXI_LCC_WVALID,
    output	wire                      S_AXI_LCC_WREADY,
    input	wire [31:0]               S_AXI_LCC_WDATA,
    input	wire [3:0]                S_AXI_LCC_WSTRB,
    output	wire                      S_AXI_LCC_BVALID,
    input	wire                      S_AXI_LCC_BREADY,
    output	wire [1:0]                S_AXI_LCC_BRESP,
    input	wire                      S_AXI_LCC_ARVALID,
    output	wire                      S_AXI_LCC_ARREADY,
    input	wire [31:0]               S_AXI_LCC_ARADDR,
    input	wire [2:0]                S_AXI_LCC_ARPROT,
    output	wire                      S_AXI_LCC_RVALID,
    input	wire                      S_AXI_LCC_RREADY,
    output	wire [31:0]               S_AXI_LCC_RDATA,
    output	wire [1:0]                S_AXI_LCC_RRESP,
    
    input wire [1:0] S_AXI_LCC_ARBURST,
    input wire [2:0] S_AXI_LCC_ARSIZE,
    input wire [7:0] S_AXI_LCC_ARLEN,
    input wire [31:0] S_AXI_LCC_ARUSER,
    input wire [18:0] S_AXI_LCC_ARID,
    input wire S_AXI_LCC_ARLOCK,
    output wire [18:0]           S_AXI_LCC_RID,
    output wire                   S_AXI_LCC_RLAST,
    input wire [             1:0] S_AXI_LCC_AWBURST,
    input wire [             2:0] S_AXI_LCC_AWSIZE,
    input wire [             7:0] S_AXI_LCC_AWLEN,
    input wire [31:0] S_AXI_LCC_AWUSER,
    input wire [18:0] S_AXI_LCC_AWID,
    input wire                    S_AXI_LCC_AWLOCK,
    input  wire                  S_AXI_LCC_WLAST,
    output wire [18:0] S_AXI_LCC_BID,

    // OTP
    input	wire                      S_AXI_OTP_AWVALID,
    output	wire                      S_AXI_OTP_AWREADY,
    input	wire [31:0]               S_AXI_OTP_AWADDR,
    input	wire [2:0]                S_AXI_OTP_AWPROT,
    input	wire                      S_AXI_OTP_WVALID,
    output	wire                      S_AXI_OTP_WREADY,
    input	wire [31:0]               S_AXI_OTP_WDATA,
    input	wire [3:0]                S_AXI_OTP_WSTRB,
    output	wire                      S_AXI_OTP_BVALID,
    input	wire                      S_AXI_OTP_BREADY,
    output	wire [1:0]                S_AXI_OTP_BRESP,
    input	wire                      S_AXI_OTP_ARVALID,
    output	wire                      S_AXI_OTP_ARREADY,
    input	wire [31:0]               S_AXI_OTP_ARADDR,
    input	wire [2:0]                S_AXI_OTP_ARPROT,
    output	wire                      S_AXI_OTP_RVALID,
    input	wire                      S_AXI_OTP_RREADY,
    output	wire [31:0]               S_AXI_OTP_RDATA,
    output	wire [1:0]                S_AXI_OTP_RRESP,
    
    input wire [1:0] S_AXI_OTP_ARBURST,
    input wire [2:0] S_AXI_OTP_ARSIZE,
    input wire [7:0] S_AXI_OTP_ARLEN,
    input wire [31:0] S_AXI_OTP_ARUSER,
    input wire [18:0] S_AXI_OTP_ARID,
    input wire S_AXI_OTP_ARLOCK,
    output wire [18:0]           S_AXI_OTP_RID,
    output wire                   S_AXI_OTP_RLAST,
    input wire [             1:0] S_AXI_OTP_AWBURST,
    input wire [             2:0] S_AXI_OTP_AWSIZE,
    input wire [             7:0] S_AXI_OTP_AWLEN,
    input wire [31:0] S_AXI_OTP_AWUSER,
    input wire [18:0] S_AXI_OTP_AWID,
    input wire                    S_AXI_OTP_AWLOCK,
    input  wire                  S_AXI_OTP_WLAST,
    output wire [18:0] S_AXI_OTP_BID,

    // ROM AXI Interface
    input  wire                       rom_backdoor_clk,
    input  wire                       rom_backdoor_en,
    input  wire [3:0]                 rom_backdoor_we,
    input  wire [16:0]                rom_backdoor_addr,
    input  wire [31:0]                rom_backdoor_din,
    output wire [31:0]                rom_backdoor_dout,
    input  wire                       rom_backdoor_rst,

    // MCU ROM Backdoor Interface
    input  wire        mcu_rom_backdoor_clk,
    input  wire        mcu_rom_backdoor_en,
    input  wire [3:0]  mcu_rom_backdoor_we,
    input  wire [31:0] mcu_rom_backdoor_addr,
    input  wire [31:0] mcu_rom_backdoor_din,
    output wire [31:0] mcu_rom_backdoor_dout,
    input  wire        mcu_rom_backdoor_rst,

    // JTAG Interface
    input wire [14:0]                  jtag_in,     // JTAG input signals concatenated
    output wire [14:0]                 jtag_out,    // JTAG tdo

    // FPGA Realtime register AXI Interface
    input	wire                      S_AXI_WRAPPER_ARESETN,
    input	wire                      S_AXI_WRAPPER_AWVALID,
    output	wire                      S_AXI_WRAPPER_AWREADY,
    input	wire [31:0]               S_AXI_WRAPPER_AWADDR,
    input	wire [2:0]                S_AXI_WRAPPER_AWPROT,
    input	wire                      S_AXI_WRAPPER_WVALID,
    output	wire                      S_AXI_WRAPPER_WREADY,
    input	wire [31:0]               S_AXI_WRAPPER_WDATA,
    input	wire [3:0]                S_AXI_WRAPPER_WSTRB,
    output	wire                      S_AXI_WRAPPER_BVALID,
    input	wire                      S_AXI_WRAPPER_BREADY,
    output	wire [1:0]                S_AXI_WRAPPER_BRESP,
    input	wire                      S_AXI_WRAPPER_ARVALID,
    output	wire                      S_AXI_WRAPPER_ARREADY,
    input	wire [31:0]               S_AXI_WRAPPER_ARADDR,
    input	wire [2:0]                S_AXI_WRAPPER_ARPROT,
    output	wire                      S_AXI_WRAPPER_RVALID,
    input	wire                      S_AXI_WRAPPER_RREADY,
    output	wire [31:0]               S_AXI_WRAPPER_RDATA,
    output	wire [1:0]                S_AXI_WRAPPER_RRESP

    // I3C
    //output SDA_UP,
    //output SDA_PUSH,
    //output SDA_PULL,
    //input  SDA,
    //output SCL_UP,
    //output SCL_PUSH,
    //output SCL_PULL,
    //input  SCL
    );

caliptra_wrapper_top cptra_wrapper (
    .core_clk(core_clk),
    .i3c_clk(i3c_clk),


    .axi_i3c_scl_t(axi_i3c_scl_t),
    .axi_i3c_scl_o(axi_i3c_scl_o),
    .axi_i3c_scl_pullup_en(axi_i3c_scl_pullup_en),
    .axi_i3c_sda_t(axi_i3c_sda_t),
    .axi_i3c_sda_o(axi_i3c_sda_o),
    .axi_i3c_sda_pullup_en(axi_i3c_sda_pullup_en),
    .SCL(SCL),
    .SDA(SDA),

    // Caliptra AXI Interface
    .S_AXI_CALIPTRA_AWADDR(S_AXI_CALIPTRA_AWADDR),
    .S_AXI_CALIPTRA_AWBURST(S_AXI_CALIPTRA_AWBURST),
    .S_AXI_CALIPTRA_AWSIZE(S_AXI_CALIPTRA_AWSIZE),
    .S_AXI_CALIPTRA_AWLEN(S_AXI_CALIPTRA_AWLEN),
    .S_AXI_CALIPTRA_AWUSER(S_AXI_CALIPTRA_AWUSER),
    .S_AXI_CALIPTRA_AWID(S_AXI_CALIPTRA_AWID),
    .S_AXI_CALIPTRA_AWLOCK(S_AXI_CALIPTRA_AWLOCK),
    .S_AXI_CALIPTRA_AWVALID(S_AXI_CALIPTRA_AWVALID),
    .S_AXI_CALIPTRA_AWREADY(S_AXI_CALIPTRA_AWREADY),
    .S_AXI_CALIPTRA_WDATA(S_AXI_CALIPTRA_WDATA),
    .S_AXI_CALIPTRA_WSTRB(S_AXI_CALIPTRA_WSTRB),
    .S_AXI_CALIPTRA_WVALID(S_AXI_CALIPTRA_WVALID),
    .S_AXI_CALIPTRA_WREADY(S_AXI_CALIPTRA_WREADY),
    .S_AXI_CALIPTRA_WLAST(S_AXI_CALIPTRA_WLAST),
    .S_AXI_CALIPTRA_BRESP(S_AXI_CALIPTRA_BRESP),
    .S_AXI_CALIPTRA_BID(S_AXI_CALIPTRA_BID),
    .S_AXI_CALIPTRA_BVALID(S_AXI_CALIPTRA_BVALID),
    .S_AXI_CALIPTRA_BREADY(S_AXI_CALIPTRA_BREADY),
    .S_AXI_CALIPTRA_ARADDR(S_AXI_CALIPTRA_ARADDR),
    .S_AXI_CALIPTRA_ARBURST(S_AXI_CALIPTRA_ARBURST),
    .S_AXI_CALIPTRA_ARSIZE(S_AXI_CALIPTRA_ARSIZE),
    .S_AXI_CALIPTRA_ARLEN(S_AXI_CALIPTRA_ARLEN),
    .S_AXI_CALIPTRA_ARUSER(S_AXI_CALIPTRA_ARUSER),
    .S_AXI_CALIPTRA_ARID(S_AXI_CALIPTRA_ARID),
    .S_AXI_CALIPTRA_ARLOCK(S_AXI_CALIPTRA_ARLOCK),
    .S_AXI_CALIPTRA_ARVALID(S_AXI_CALIPTRA_ARVALID),
    .S_AXI_CALIPTRA_ARREADY(S_AXI_CALIPTRA_ARREADY),
    .S_AXI_CALIPTRA_RDATA(S_AXI_CALIPTRA_RDATA),
    .S_AXI_CALIPTRA_RRESP(S_AXI_CALIPTRA_RRESP),
    .S_AXI_CALIPTRA_RID(S_AXI_CALIPTRA_RID),
    .S_AXI_CALIPTRA_RLAST(S_AXI_CALIPTRA_RLAST),
    .S_AXI_CALIPTRA_RVALID(S_AXI_CALIPTRA_RVALID),
    .S_AXI_CALIPTRA_RREADY(S_AXI_CALIPTRA_RREADY),

    // Caliptra M_AXI Interface
    .M_AXI_CALIPTRA_AWADDR(M_AXI_CALIPTRA_AWADDR),
    .M_AXI_CALIPTRA_AWBURST(M_AXI_CALIPTRA_AWBURST),
    .M_AXI_CALIPTRA_AWSIZE(M_AXI_CALIPTRA_AWSIZE),
    .M_AXI_CALIPTRA_AWLEN(M_AXI_CALIPTRA_AWLEN),
    .M_AXI_CALIPTRA_AWUSER(M_AXI_CALIPTRA_AWUSER),
    .M_AXI_CALIPTRA_AWID(M_AXI_CALIPTRA_AWID),
    .M_AXI_CALIPTRA_AWLOCK(M_AXI_CALIPTRA_AWLOCK),
    .M_AXI_CALIPTRA_AWVALID(M_AXI_CALIPTRA_AWVALID),
    .M_AXI_CALIPTRA_AWREADY(M_AXI_CALIPTRA_AWREADY),
    // W
    .M_AXI_CALIPTRA_WDATA(M_AXI_CALIPTRA_WDATA),
    .M_AXI_CALIPTRA_WSTRB(M_AXI_CALIPTRA_WSTRB),
    .M_AXI_CALIPTRA_WVALID(M_AXI_CALIPTRA_WVALID),
    .M_AXI_CALIPTRA_WREADY(M_AXI_CALIPTRA_WREADY),
    .M_AXI_CALIPTRA_WLAST(M_AXI_CALIPTRA_WLAST),
    // B
    .M_AXI_CALIPTRA_BRESP(M_AXI_CALIPTRA_BRESP),
    .M_AXI_CALIPTRA_BID(M_AXI_CALIPTRA_BID),
    .M_AXI_CALIPTRA_BVALID(M_AXI_CALIPTRA_BVALID),
    .M_AXI_CALIPTRA_BREADY(M_AXI_CALIPTRA_BREADY),
    // AR
    .M_AXI_CALIPTRA_ARADDR(M_AXI_CALIPTRA_ARADDR),
    .M_AXI_CALIPTRA_ARBURST(M_AXI_CALIPTRA_ARBURST),
    .M_AXI_CALIPTRA_ARSIZE(M_AXI_CALIPTRA_ARSIZE),
    .M_AXI_CALIPTRA_ARLEN(M_AXI_CALIPTRA_ARLEN),
    .M_AXI_CALIPTRA_ARUSER(M_AXI_CALIPTRA_ARUSER),
    .M_AXI_CALIPTRA_ARID(M_AXI_CALIPTRA_ARID),
    .M_AXI_CALIPTRA_ARLOCK(M_AXI_CALIPTRA_ARLOCK),
    .M_AXI_CALIPTRA_ARVALID(M_AXI_CALIPTRA_ARVALID),
    .M_AXI_CALIPTRA_ARREADY(M_AXI_CALIPTRA_ARREADY),
    // R
    .M_AXI_CALIPTRA_RDATA(M_AXI_CALIPTRA_RDATA),
    .M_AXI_CALIPTRA_RRESP(M_AXI_CALIPTRA_RRESP),
    .M_AXI_CALIPTRA_RID(M_AXI_CALIPTRA_RID),
    .M_AXI_CALIPTRA_RLAST(M_AXI_CALIPTRA_RLAST),
    .M_AXI_CALIPTRA_RVALID(M_AXI_CALIPTRA_RVALID),
    .M_AXI_CALIPTRA_RREADY(M_AXI_CALIPTRA_RREADY),


    // MCI AXI Interface
    .S_AXI_MCI_AWADDR(S_AXI_MCI_AWADDR),
    .S_AXI_MCI_AWBURST(S_AXI_MCI_AWBURST),
    .S_AXI_MCI_AWSIZE(S_AXI_MCI_AWSIZE),
    .S_AXI_MCI_AWLEN(S_AXI_MCI_AWLEN),
    .S_AXI_MCI_AWUSER(S_AXI_MCI_AWUSER),
    .S_AXI_MCI_AWID(S_AXI_MCI_AWID),
    .S_AXI_MCI_AWLOCK(S_AXI_MCI_AWLOCK),
    .S_AXI_MCI_AWVALID(S_AXI_MCI_AWVALID),
    .S_AXI_MCI_AWREADY(S_AXI_MCI_AWREADY),
    .S_AXI_MCI_WDATA(S_AXI_MCI_WDATA),
    .S_AXI_MCI_WSTRB(S_AXI_MCI_WSTRB),
    .S_AXI_MCI_WVALID(S_AXI_MCI_WVALID),
    .S_AXI_MCI_WREADY(S_AXI_MCI_WREADY),
    .S_AXI_MCI_WLAST(S_AXI_MCI_WLAST),
    .S_AXI_MCI_BRESP(S_AXI_MCI_BRESP),
    .S_AXI_MCI_BID(S_AXI_MCI_BID),
    .S_AXI_MCI_BVALID(S_AXI_MCI_BVALID),
    .S_AXI_MCI_BREADY(S_AXI_MCI_BREADY),
    .S_AXI_MCI_ARADDR(S_AXI_MCI_ARADDR),
    .S_AXI_MCI_ARBURST(S_AXI_MCI_ARBURST),
    .S_AXI_MCI_ARSIZE(S_AXI_MCI_ARSIZE),
    .S_AXI_MCI_ARLEN(S_AXI_MCI_ARLEN),
    .S_AXI_MCI_ARUSER(S_AXI_MCI_ARUSER),
    .S_AXI_MCI_ARID(S_AXI_MCI_ARID),
    .S_AXI_MCI_ARLOCK(S_AXI_MCI_ARLOCK),
    .S_AXI_MCI_ARVALID(S_AXI_MCI_ARVALID),
    .S_AXI_MCI_ARREADY(S_AXI_MCI_ARREADY),
    .S_AXI_MCI_RDATA(S_AXI_MCI_RDATA),
    .S_AXI_MCI_RRESP(S_AXI_MCI_RRESP),
    .S_AXI_MCI_RID(S_AXI_MCI_RID),
    .S_AXI_MCI_RLAST(S_AXI_MCI_RLAST),
    .S_AXI_MCI_RVALID(S_AXI_MCI_RVALID),
    .S_AXI_MCI_RREADY(S_AXI_MCI_RREADY),

    // MCI ROM AXI Interface
    .S_AXI_MCU_ROM_AWADDR(S_AXI_MCU_ROM_AWADDR),
    .S_AXI_MCU_ROM_AWBURST(S_AXI_MCU_ROM_AWBURST),
    .S_AXI_MCU_ROM_AWSIZE(S_AXI_MCU_ROM_AWSIZE),
    .S_AXI_MCU_ROM_AWLEN(S_AXI_MCU_ROM_AWLEN),
    .S_AXI_MCU_ROM_AWUSER(S_AXI_MCU_ROM_AWUSER),
    .S_AXI_MCU_ROM_AWID(S_AXI_MCU_ROM_AWID),
    .S_AXI_MCU_ROM_AWLOCK(S_AXI_MCU_ROM_AWLOCK),
    .S_AXI_MCU_ROM_AWVALID(S_AXI_MCU_ROM_AWVALID),
    .S_AXI_MCU_ROM_AWREADY(S_AXI_MCU_ROM_AWREADY),
    .S_AXI_MCU_ROM_WDATA(S_AXI_MCU_ROM_WDATA),
    .S_AXI_MCU_ROM_WSTRB(S_AXI_MCU_ROM_WSTRB),
    .S_AXI_MCU_ROM_WVALID(S_AXI_MCU_ROM_WVALID),
    .S_AXI_MCU_ROM_WREADY(S_AXI_MCU_ROM_WREADY),
    .S_AXI_MCU_ROM_WLAST(S_AXI_MCU_ROM_WLAST),
    .S_AXI_MCU_ROM_BRESP(S_AXI_MCU_ROM_BRESP),
    .S_AXI_MCU_ROM_BID(S_AXI_MCU_ROM_BID),
    .S_AXI_MCU_ROM_BVALID(S_AXI_MCU_ROM_BVALID),
    .S_AXI_MCU_ROM_BREADY(S_AXI_MCU_ROM_BREADY),
    .S_AXI_MCU_ROM_ARADDR(S_AXI_MCU_ROM_ARADDR),
    .S_AXI_MCU_ROM_ARBURST(S_AXI_MCU_ROM_ARBURST),
    .S_AXI_MCU_ROM_ARSIZE(S_AXI_MCU_ROM_ARSIZE),
    .S_AXI_MCU_ROM_ARLEN(S_AXI_MCU_ROM_ARLEN),
    .S_AXI_MCU_ROM_ARUSER(S_AXI_MCU_ROM_ARUSER),
    .S_AXI_MCU_ROM_ARID(S_AXI_MCU_ROM_ARID),
    .S_AXI_MCU_ROM_ARLOCK(S_AXI_MCU_ROM_ARLOCK),
    .S_AXI_MCU_ROM_ARVALID(S_AXI_MCU_ROM_ARVALID),
    .S_AXI_MCU_ROM_ARREADY(S_AXI_MCU_ROM_ARREADY),
    .S_AXI_MCU_ROM_RDATA(S_AXI_MCU_ROM_RDATA),
    .S_AXI_MCU_ROM_RRESP(S_AXI_MCU_ROM_RRESP),
    .S_AXI_MCU_ROM_RID(S_AXI_MCU_ROM_RID),
    .S_AXI_MCU_ROM_RLAST(S_AXI_MCU_ROM_RLAST),
    .S_AXI_MCU_ROM_RVALID(S_AXI_MCU_ROM_RVALID),
    .S_AXI_MCU_ROM_RREADY(S_AXI_MCU_ROM_RREADY),

    // Caliptra M_AXI Interface
    .M_AXI_MCI_AWADDR(M_AXI_MCI_AWADDR),
    .M_AXI_MCI_AWBURST(M_AXI_MCI_AWBURST),
    .M_AXI_MCI_AWSIZE(M_AXI_MCI_AWSIZE),
    .M_AXI_MCI_AWLEN(M_AXI_MCI_AWLEN),
    .M_AXI_MCI_AWUSER(M_AXI_MCI_AWUSER),
    .M_AXI_MCI_AWID(M_AXI_MCI_AWID),
    .M_AXI_MCI_AWLOCK(M_AXI_MCI_AWLOCK),
    .M_AXI_MCI_AWVALID(M_AXI_MCI_AWVALID),
    .M_AXI_MCI_AWREADY(M_AXI_MCI_AWREADY),
    // W
    .M_AXI_MCI_WDATA(M_AXI_MCI_WDATA),
    .M_AXI_MCI_WSTRB(M_AXI_MCI_WSTRB),
    .M_AXI_MCI_WVALID(M_AXI_MCI_WVALID),
    .M_AXI_MCI_WREADY(M_AXI_MCI_WREADY),
    .M_AXI_MCI_WLAST(M_AXI_MCI_WLAST),
    // B
    .M_AXI_MCI_BRESP(M_AXI_MCI_BRESP),
    .M_AXI_MCI_BID(M_AXI_MCI_BID),
    .M_AXI_MCI_BVALID(M_AXI_MCI_BVALID),
    .M_AXI_MCI_BREADY(M_AXI_MCI_BREADY),
    // AR
    .M_AXI_MCI_ARADDR(M_AXI_MCI_ARADDR),
    .M_AXI_MCI_ARBURST(M_AXI_MCI_ARBURST),
    .M_AXI_MCI_ARSIZE(M_AXI_MCI_ARSIZE),
    .M_AXI_MCI_ARLEN(M_AXI_MCI_ARLEN),
    .M_AXI_MCI_ARUSER(M_AXI_MCI_ARUSER),
    .M_AXI_MCI_ARID(M_AXI_MCI_ARID),
    .M_AXI_MCI_ARLOCK(M_AXI_MCI_ARLOCK),
    .M_AXI_MCI_ARVALID(M_AXI_MCI_ARVALID),
    .M_AXI_MCI_ARREADY(M_AXI_MCI_ARREADY),
    // R
    .M_AXI_MCI_RDATA(M_AXI_MCI_RDATA),
    .M_AXI_MCI_RRESP(M_AXI_MCI_RRESP),
    .M_AXI_MCI_RID(M_AXI_MCI_RID),
    .M_AXI_MCI_RLAST(M_AXI_MCI_RLAST),
    .M_AXI_MCI_RVALID(M_AXI_MCI_RVALID),
    .M_AXI_MCI_RREADY(M_AXI_MCI_RREADY),

    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_LSU_AWVALID(M_AXI_MCU_LSU_AWVALID),
    .M_AXI_MCU_LSU_AWREADY(M_AXI_MCU_LSU_AWREADY),
    .M_AXI_MCU_LSU_AWID(M_AXI_MCU_LSU_AWID),
    .M_AXI_MCU_LSU_AWADDR(M_AXI_MCU_LSU_AWADDR),
    .M_AXI_MCU_LSU_AWREGION(M_AXI_MCU_LSU_AWREGION),
    .M_AXI_MCU_LSU_AWLEN(M_AXI_MCU_LSU_AWLEN),
    .M_AXI_MCU_LSU_AWSIZE(M_AXI_MCU_LSU_AWSIZE),
    .M_AXI_MCU_LSU_AWBURST(M_AXI_MCU_LSU_AWBURST),
    .M_AXI_MCU_LSU_AWLOCK(M_AXI_MCU_LSU_AWLOCK),
    .M_AXI_MCU_LSU_AWCACHE(M_AXI_MCU_LSU_AWCACHE),
    .M_AXI_MCU_LSU_AWPROT(M_AXI_MCU_LSU_AWPROT),
    .M_AXI_MCU_LSU_AWQOS(M_AXI_MCU_LSU_AWQOS),

    .M_AXI_MCU_LSU_WVALID(M_AXI_MCU_LSU_WVALID),
    .M_AXI_MCU_LSU_WREADY(M_AXI_MCU_LSU_WREADY),
    .M_AXI_MCU_LSU_WDATA(M_AXI_MCU_LSU_WDATA),
    .M_AXI_MCU_LSU_WSTRB(M_AXI_MCU_LSU_WSTRB),
    .M_AXI_MCU_LSU_WLAST(M_AXI_MCU_LSU_WLAST),

    .M_AXI_MCU_LSU_BVALID(M_AXI_MCU_LSU_BVALID),
    .M_AXI_MCU_LSU_BREADY(M_AXI_MCU_LSU_BREADY),
    .M_AXI_MCU_LSU_BRESP(M_AXI_MCU_LSU_BRESP),
    .M_AXI_MCU_LSU_BID(M_AXI_MCU_LSU_BID),

    // AXI Read Channels
    .M_AXI_MCU_LSU_ARVALID(M_AXI_MCU_LSU_ARVALID),
    .M_AXI_MCU_LSU_ARREADY(M_AXI_MCU_LSU_ARREADY),
    .M_AXI_MCU_LSU_ARID(M_AXI_MCU_LSU_ARID),
    .M_AXI_MCU_LSU_ARADDR(M_AXI_MCU_LSU_ARADDR),
    .M_AXI_MCU_LSU_ARREGION(M_AXI_MCU_LSU_ARREGION),
    .M_AXI_MCU_LSU_ARLEN(M_AXI_MCU_LSU_ARLEN),
    .M_AXI_MCU_LSU_ARSIZE(M_AXI_MCU_LSU_ARSIZE),
    .M_AXI_MCU_LSU_ARBURST(M_AXI_MCU_LSU_ARBURST),
    .M_AXI_MCU_LSU_ARLOCK(M_AXI_MCU_LSU_ARLOCK),
    .M_AXI_MCU_LSU_ARCACHE(M_AXI_MCU_LSU_ARCACHE),
    .M_AXI_MCU_LSU_ARPROT(M_AXI_MCU_LSU_ARPROT),
    .M_AXI_MCU_LSU_ARQOS(M_AXI_MCU_LSU_ARQOS),

    .M_AXI_MCU_LSU_RVALID(M_AXI_MCU_LSU_RVALID),
    .M_AXI_MCU_LSU_RREADY(M_AXI_MCU_LSU_RREADY),
    .M_AXI_MCU_LSU_RID(M_AXI_MCU_LSU_RID),
    .M_AXI_MCU_LSU_RDATA(M_AXI_MCU_LSU_RDATA),
    .M_AXI_MCU_LSU_RRESP(M_AXI_MCU_LSU_RRESP),
    .M_AXI_MCU_LSU_RLAST(M_AXI_MCU_LSU_RLAST),

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_IFU_AWVALID(M_AXI_MCU_IFU_AWVALID),
    .M_AXI_MCU_IFU_AWREADY(M_AXI_MCU_IFU_AWREADY),
    .M_AXI_MCU_IFU_AWID(M_AXI_MCU_IFU_AWID),
    .M_AXI_MCU_IFU_AWADDR(M_AXI_MCU_IFU_AWADDR),
    .M_AXI_MCU_IFU_AWREGION(M_AXI_MCU_IFU_AWREGION),
    .M_AXI_MCU_IFU_AWLEN(M_AXI_MCU_IFU_AWLEN),
    .M_AXI_MCU_IFU_AWSIZE(M_AXI_MCU_IFU_AWSIZE),
    .M_AXI_MCU_IFU_AWBURST(M_AXI_MCU_IFU_AWBURST),
    .M_AXI_MCU_IFU_AWLOCK(M_AXI_MCU_IFU_AWLOCK),
    .M_AXI_MCU_IFU_AWCACHE(M_AXI_MCU_IFU_AWCACHE),
    .M_AXI_MCU_IFU_AWPROT(M_AXI_MCU_IFU_AWPROT),
    .M_AXI_MCU_IFU_AWQOS(M_AXI_MCU_IFU_AWQOS),

    .M_AXI_MCU_IFU_WVALID(M_AXI_MCU_IFU_WVALID),
    .M_AXI_MCU_IFU_WREADY(M_AXI_MCU_IFU_WREADY),
    .M_AXI_MCU_IFU_WDATA(M_AXI_MCU_IFU_WDATA),
    .M_AXI_MCU_IFU_WSTRB(M_AXI_MCU_IFU_WSTRB),
    .M_AXI_MCU_IFU_WLAST(M_AXI_MCU_IFU_WLAST),

    .M_AXI_MCU_IFU_BVALID(M_AXI_MCU_IFU_BVALID),
    .M_AXI_MCU_IFU_BREADY(M_AXI_MCU_IFU_BREADY),
    .M_AXI_MCU_IFU_BRESP(M_AXI_MCU_IFU_BRESP),
    .M_AXI_MCU_IFU_BID(M_AXI_MCU_IFU_BID),

    // AXI Read Channels
    .M_AXI_MCU_IFU_ARVALID(M_AXI_MCU_IFU_ARVALID),
    .M_AXI_MCU_IFU_ARREADY(M_AXI_MCU_IFU_ARREADY),
    .M_AXI_MCU_IFU_ARID(M_AXI_MCU_IFU_ARID),
    .M_AXI_MCU_IFU_ARADDR(M_AXI_MCU_IFU_ARADDR),
    .M_AXI_MCU_IFU_ARREGION(M_AXI_MCU_IFU_ARREGION),
    .M_AXI_MCU_IFU_ARLEN(M_AXI_MCU_IFU_ARLEN),
    .M_AXI_MCU_IFU_ARSIZE(M_AXI_MCU_IFU_ARSIZE),
    .M_AXI_MCU_IFU_ARBURST(M_AXI_MCU_IFU_ARBURST),
    .M_AXI_MCU_IFU_ARLOCK(M_AXI_MCU_IFU_ARLOCK),
    .M_AXI_MCU_IFU_ARCACHE(M_AXI_MCU_IFU_ARCACHE),
    .M_AXI_MCU_IFU_ARPROT(M_AXI_MCU_IFU_ARPROT),
    .M_AXI_MCU_IFU_ARQOS(M_AXI_MCU_IFU_ARQOS),

    .M_AXI_MCU_IFU_RVALID(M_AXI_MCU_IFU_RVALID),
    .M_AXI_MCU_IFU_RREADY(M_AXI_MCU_IFU_RREADY),
    .M_AXI_MCU_IFU_RID(M_AXI_MCU_IFU_RID),
    .M_AXI_MCU_IFU_RDATA(M_AXI_MCU_IFU_RDATA),
    .M_AXI_MCU_IFU_RRESP(M_AXI_MCU_IFU_RRESP),
    .M_AXI_MCU_IFU_RLAST(M_AXI_MCU_IFU_RLAST),

    //-------------------------- MCU SB AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_SB_AWVALID(M_AXI_MCU_SB_AWVALID),
    .M_AXI_MCU_SB_AWREADY(M_AXI_MCU_SB_AWREADY),
    .M_AXI_MCU_SB_AWID(M_AXI_MCU_SB_AWID),
    .M_AXI_MCU_SB_AWADDR(M_AXI_MCU_SB_AWADDR),
    .M_AXI_MCU_SB_AWREGION(M_AXI_MCU_SB_AWREGION),
    .M_AXI_MCU_SB_AWLEN(M_AXI_MCU_SB_AWLEN),
    .M_AXI_MCU_SB_AWSIZE(M_AXI_MCU_SB_AWSIZE),
    .M_AXI_MCU_SB_AWBURST(M_AXI_MCU_SB_AWBURST),
    .M_AXI_MCU_SB_AWLOCK(M_AXI_MCU_SB_AWLOCK),
    .M_AXI_MCU_SB_AWCACHE(M_AXI_MCU_SB_AWCACHE),
    .M_AXI_MCU_SB_AWPROT(M_AXI_MCU_SB_AWPROT),
    .M_AXI_MCU_SB_AWQOS(M_AXI_MCU_SB_AWQOS),

    .M_AXI_MCU_SB_WVALID(M_AXI_MCU_SB_WVALID),
    .M_AXI_MCU_SB_WREADY(M_AXI_MCU_SB_WREADY),
    .M_AXI_MCU_SB_WDATA(M_AXI_MCU_SB_WDATA),
    .M_AXI_MCU_SB_WSTRB(M_AXI_MCU_SB_WSTRB),
    .M_AXI_MCU_SB_WLAST(M_AXI_MCU_SB_WLAST),

    .M_AXI_MCU_SB_BVALID(M_AXI_MCU_SB_BVALID),
    .M_AXI_MCU_SB_BREADY(M_AXI_MCU_SB_BREADY),
    .M_AXI_MCU_SB_BRESP(M_AXI_MCU_SB_BRESP),
    .M_AXI_MCU_SB_BID(M_AXI_MCU_SB_BID),

    // AXI Read Channels
    .M_AXI_MCU_SB_ARVALID(M_AXI_MCU_SB_ARVALID),
    .M_AXI_MCU_SB_ARREADY(M_AXI_MCU_SB_ARREADY),
    .M_AXI_MCU_SB_ARID(M_AXI_MCU_SB_ARID),
    .M_AXI_MCU_SB_ARADDR(M_AXI_MCU_SB_ARADDR),
    .M_AXI_MCU_SB_ARREGION(M_AXI_MCU_SB_ARREGION),
    .M_AXI_MCU_SB_ARLEN(M_AXI_MCU_SB_ARLEN),
    .M_AXI_MCU_SB_ARSIZE(M_AXI_MCU_SB_ARSIZE),
    .M_AXI_MCU_SB_ARBURST(M_AXI_MCU_SB_ARBURST),
    .M_AXI_MCU_SB_ARLOCK(M_AXI_MCU_SB_ARLOCK),
    .M_AXI_MCU_SB_ARCACHE(M_AXI_MCU_SB_ARCACHE),
    .M_AXI_MCU_SB_ARPROT(M_AXI_MCU_SB_ARPROT),
    .M_AXI_MCU_SB_ARQOS(M_AXI_MCU_SB_ARQOS),

    .M_AXI_MCU_SB_RVALID(M_AXI_MCU_SB_RVALID),
    .M_AXI_MCU_SB_RREADY(M_AXI_MCU_SB_RREADY),
    .M_AXI_MCU_SB_RID(M_AXI_MCU_SB_RID),
    .M_AXI_MCU_SB_RDATA(M_AXI_MCU_SB_RDATA),
    .M_AXI_MCU_SB_RRESP(M_AXI_MCU_SB_RRESP),
    .M_AXI_MCU_SB_RLAST(M_AXI_MCU_SB_RLAST),

    // I3C
    .S_AXI_I3C_AWVALID(S_AXI_I3C_AWVALID),
    .S_AXI_I3C_AWREADY(S_AXI_I3C_AWREADY),
    .S_AXI_I3C_AWADDR(S_AXI_I3C_AWADDR),
    .S_AXI_I3C_AWPROT(S_AXI_I3C_AWPROT),
    .S_AXI_I3C_WVALID(S_AXI_I3C_WVALID),
    .S_AXI_I3C_WREADY(S_AXI_I3C_WREADY),
    .S_AXI_I3C_WDATA(S_AXI_I3C_WDATA),
    .S_AXI_I3C_WSTRB(S_AXI_I3C_WSTRB),
    .S_AXI_I3C_BVALID(S_AXI_I3C_BVALID),
    .S_AXI_I3C_BREADY(S_AXI_I3C_BREADY),
    .S_AXI_I3C_BRESP(S_AXI_I3C_BRESP),
    .S_AXI_I3C_ARVALID(S_AXI_I3C_ARVALID),
    .S_AXI_I3C_ARREADY(S_AXI_I3C_ARREADY),
    .S_AXI_I3C_ARADDR(S_AXI_I3C_ARADDR),
    .S_AXI_I3C_ARPROT(S_AXI_I3C_ARPROT),
    .S_AXI_I3C_RVALID(S_AXI_I3C_RVALID),
    .S_AXI_I3C_RREADY(S_AXI_I3C_RREADY),
    .S_AXI_I3C_RDATA(S_AXI_I3C_RDATA),
    .S_AXI_I3C_RRESP(S_AXI_I3C_RRESP),
    .S_AXI_I3C_ARBURST(S_AXI_I3C_ARBURST),
    .S_AXI_I3C_ARSIZE(S_AXI_I3C_ARSIZE),
    .S_AXI_I3C_ARLEN(S_AXI_I3C_ARLEN),
    .S_AXI_I3C_ARUSER(S_AXI_I3C_ARUSER),
    .S_AXI_I3C_ARID(S_AXI_I3C_ARID),
    .S_AXI_I3C_ARLOCK(S_AXI_I3C_ARLOCK),
    .S_AXI_I3C_RID(S_AXI_I3C_RID),
    .S_AXI_I3C_RLAST(S_AXI_I3C_RLAST),
    .S_AXI_I3C_AWBURST(S_AXI_I3C_AWBURST),
    .S_AXI_I3C_AWSIZE(S_AXI_I3C_AWSIZE),
    .S_AXI_I3C_AWLEN(S_AXI_I3C_AWLEN),
    .S_AXI_I3C_AWUSER(S_AXI_I3C_AWUSER),
    .S_AXI_I3C_AWID(S_AXI_I3C_AWID),
    .S_AXI_I3C_AWLOCK(S_AXI_I3C_AWLOCK),
    .S_AXI_I3C_WLAST(S_AXI_I3C_WLAST),
    .S_AXI_I3C_BID(S_AXI_I3C_BID),

    // LCC
    .S_AXI_LCC_AWVALID(S_AXI_LCC_AWVALID),
    .S_AXI_LCC_AWREADY(S_AXI_LCC_AWREADY),
    .S_AXI_LCC_AWADDR(S_AXI_LCC_AWADDR),
    .S_AXI_LCC_AWPROT(S_AXI_LCC_AWPROT),
    .S_AXI_LCC_WVALID(S_AXI_LCC_WVALID),
    .S_AXI_LCC_WREADY(S_AXI_LCC_WREADY),
    .S_AXI_LCC_WDATA(S_AXI_LCC_WDATA),
    .S_AXI_LCC_WSTRB(S_AXI_LCC_WSTRB),
    .S_AXI_LCC_BVALID(S_AXI_LCC_BVALID),
    .S_AXI_LCC_BREADY(S_AXI_LCC_BREADY),
    .S_AXI_LCC_BRESP(S_AXI_LCC_BRESP),
    .S_AXI_LCC_ARVALID(S_AXI_LCC_ARVALID),
    .S_AXI_LCC_ARREADY(S_AXI_LCC_ARREADY),
    .S_AXI_LCC_ARADDR(S_AXI_LCC_ARADDR),
    .S_AXI_LCC_ARPROT(S_AXI_LCC_ARPROT),
    .S_AXI_LCC_RVALID(S_AXI_LCC_RVALID),
    .S_AXI_LCC_RREADY(S_AXI_LCC_RREADY),
    .S_AXI_LCC_RDATA(S_AXI_LCC_RDATA),
    .S_AXI_LCC_RRESP(S_AXI_LCC_RRESP),
    
    .S_AXI_LCC_ARBURST(S_AXI_LCC_ARBURST),
    .S_AXI_LCC_ARSIZE(S_AXI_LCC_ARSIZE),
    .S_AXI_LCC_ARLEN(S_AXI_LCC_ARLEN),
    .S_AXI_LCC_ARUSER(S_AXI_LCC_ARUSER),
    .S_AXI_LCC_ARID(S_AXI_LCC_ARID),
    .S_AXI_LCC_ARLOCK(S_AXI_LCC_ARLOCK),
    .S_AXI_LCC_RID(S_AXI_LCC_RID),
    .S_AXI_LCC_RLAST(S_AXI_LCC_RLAST),
    .S_AXI_LCC_AWBURST(S_AXI_LCC_AWBURST),
    .S_AXI_LCC_AWSIZE(S_AXI_LCC_AWSIZE),
    .S_AXI_LCC_AWLEN(S_AXI_LCC_AWLEN),
    .S_AXI_LCC_AWUSER(S_AXI_LCC_AWUSER),
    .S_AXI_LCC_AWID(S_AXI_LCC_AWID),
    .S_AXI_LCC_AWLOCK(S_AXI_LCC_AWLOCK),
    .S_AXI_LCC_WLAST(S_AXI_LCC_WLAST),
    .S_AXI_LCC_BID(S_AXI_LCC_BID),

    // OTP
    .S_AXI_OTP_AWVALID(S_AXI_OTP_AWVALID),
    .S_AXI_OTP_AWREADY(S_AXI_OTP_AWREADY),
    .S_AXI_OTP_AWADDR(S_AXI_OTP_AWADDR),
    .S_AXI_OTP_AWPROT(S_AXI_OTP_AWPROT),
    .S_AXI_OTP_WVALID(S_AXI_OTP_WVALID),
    .S_AXI_OTP_WREADY(S_AXI_OTP_WREADY),
    .S_AXI_OTP_WDATA(S_AXI_OTP_WDATA),
    .S_AXI_OTP_WSTRB(S_AXI_OTP_WSTRB),
    .S_AXI_OTP_BVALID(S_AXI_OTP_BVALID),
    .S_AXI_OTP_BREADY(S_AXI_OTP_BREADY),
    .S_AXI_OTP_BRESP(S_AXI_OTP_BRESP),
    .S_AXI_OTP_ARVALID(S_AXI_OTP_ARVALID),
    .S_AXI_OTP_ARREADY(S_AXI_OTP_ARREADY),
    .S_AXI_OTP_ARADDR(S_AXI_OTP_ARADDR),
    .S_AXI_OTP_ARPROT(S_AXI_OTP_ARPROT),
    .S_AXI_OTP_RVALID(S_AXI_OTP_RVALID),
    .S_AXI_OTP_RREADY(S_AXI_OTP_RREADY),
    .S_AXI_OTP_RDATA(S_AXI_OTP_RDATA),
    .S_AXI_OTP_RRESP(S_AXI_OTP_RRESP),
    
    .S_AXI_OTP_ARBURST(S_AXI_OTP_ARBURST),
    .S_AXI_OTP_ARSIZE(S_AXI_OTP_ARSIZE),
    .S_AXI_OTP_ARLEN(S_AXI_OTP_ARLEN),
    .S_AXI_OTP_ARUSER(S_AXI_OTP_ARUSER),
    .S_AXI_OTP_ARID(S_AXI_OTP_ARID),
    .S_AXI_OTP_ARLOCK(S_AXI_OTP_ARLOCK),
    .S_AXI_OTP_RID(S_AXI_OTP_RID),
    .S_AXI_OTP_RLAST(S_AXI_OTP_RLAST),
    .S_AXI_OTP_AWBURST(S_AXI_OTP_AWBURST),
    .S_AXI_OTP_AWSIZE(S_AXI_OTP_AWSIZE),
    .S_AXI_OTP_AWLEN(S_AXI_OTP_AWLEN),
    .S_AXI_OTP_AWUSER(S_AXI_OTP_AWUSER),
    .S_AXI_OTP_AWID(S_AXI_OTP_AWID),
    .S_AXI_OTP_AWLOCK(S_AXI_OTP_AWLOCK),
    .S_AXI_OTP_WLAST(S_AXI_OTP_WLAST),
    .S_AXI_OTP_BID(S_AXI_OTP_BID),

    // SOC access to program ROM
    .rom_backdoor_clk(rom_backdoor_clk),
    .rom_backdoor_en(rom_backdoor_en),
    .rom_backdoor_we(rom_backdoor_we),
    .rom_backdoor_addr(rom_backdoor_addr[16:2]),
    .rom_backdoor_wrdata(rom_backdoor_din),
    .rom_backdoor_rddata(rom_backdoor_dout),
    .rom_backdoor_rst(rom_backdoor_rst),

    // SOC access to program MCU ROM
    .mcu_rom_backdoor_clk(mcu_rom_backdoor_clk),
    .mcu_rom_backdoor_en(mcu_rom_backdoor_en),
    .mcu_rom_backdoor_we(mcu_rom_backdoor_we),
    .mcu_rom_backdoor_addr(mcu_rom_backdoor_addr[31:2]),
    .mcu_rom_backdoor_din(mcu_rom_backdoor_din),
    .mcu_rom_backdoor_dout(mcu_rom_backdoor_dout),
    .mcu_rom_backdoor_rst(mcu_rom_backdoor_rst),

    // EL2 JTAG interface
    .jtag_tck(jtag_in[0]),
    .jtag_tdi(jtag_in[1]),
    .jtag_tms(jtag_in[2]),
    .jtag_trst_n(jtag_in[3]),
    .jtag_tdo(jtag_out[4]),

    // MCU
    .mcu_jtag_tck_i(jtag_in[5]),
    .mcu_jtag_tms_i(jtag_in[6]),
    .mcu_jtag_tdi_i(jtag_in[7]),
    .mcu_jtag_trst_n_i(jtag_in[8]),
    .mcu_jtag_tdo_o(jtag_out[9]),
    
    .lc_jtag_tck_i(jtag_in[10]),
    .lc_jtag_tms_i(jtag_in[11]),
    .lc_jtag_tdi_i(jtag_in[12]),
    .lc_jtag_trst_n_i(jtag_in[13]),
    .lc_jtag_tdo_o(jtag_out[14]),

    // FPGA Realtime register AXI Interface
    .S_AXI_WRAPPER_ARESETN(S_AXI_WRAPPER_ARESETN),
    .S_AXI_WRAPPER_AWVALID(S_AXI_WRAPPER_AWVALID),
    .S_AXI_WRAPPER_AWREADY(S_AXI_WRAPPER_AWREADY),
    .S_AXI_WRAPPER_AWADDR(S_AXI_WRAPPER_AWADDR),
    .S_AXI_WRAPPER_AWPROT(S_AXI_WRAPPER_AWPROT),
    .S_AXI_WRAPPER_WVALID(S_AXI_WRAPPER_WVALID),
    .S_AXI_WRAPPER_WREADY(S_AXI_WRAPPER_WREADY),
    .S_AXI_WRAPPER_WDATA(S_AXI_WRAPPER_WDATA),
    .S_AXI_WRAPPER_WSTRB(S_AXI_WRAPPER_WSTRB),
    .S_AXI_WRAPPER_BVALID(S_AXI_WRAPPER_BVALID),
    .S_AXI_WRAPPER_BREADY(S_AXI_WRAPPER_BREADY),
    .S_AXI_WRAPPER_BRESP(S_AXI_WRAPPER_BRESP),
    .S_AXI_WRAPPER_ARVALID(S_AXI_WRAPPER_ARVALID),
    .S_AXI_WRAPPER_ARREADY(S_AXI_WRAPPER_ARREADY),
    .S_AXI_WRAPPER_ARADDR(S_AXI_WRAPPER_ARADDR),
    .S_AXI_WRAPPER_ARPROT(S_AXI_WRAPPER_ARPROT),
    .S_AXI_WRAPPER_RVALID(S_AXI_WRAPPER_RVALID),
    .S_AXI_WRAPPER_RREADY(S_AXI_WRAPPER_RREADY),
    .S_AXI_WRAPPER_RDATA(S_AXI_WRAPPER_RDATA),
    .S_AXI_WRAPPER_RRESP(S_AXI_WRAPPER_RRESP)

    //.SDA_UP(SDA_UP),
    //.SDA_PUSH(SDA_PUSH),
    //.SDA_PULL(SDA_PULL),
    //.SDA(SDA),
    //.SCL_UP(SCL_UP),
    //.SCL_PUSH(SCL_PUSH),
    //.SCL_PULL(SCL_PULL),
    //.SCL(SCL)
);
endmodule
