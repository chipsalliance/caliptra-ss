// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module mci_boot_seqr #(
    parameter myparam = "fixme"
) (
    input logic clk,
    input logic rst_n,

    output logic fabric_rst_b,
    output logic fc_rst_b,
    output logic lcc_rst_b,
    output logic tap_rst_b,
    output logic mcu_rst_b,
    output logic cptra_rst_b
);

endmodule
