
module caliptra_ss_package_top (
    input wire core_clk,

    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_LSU_AWVALID,
    input  wire                      M_AXI_MCU_LSU_AWREADY,
    output wire [18:0]               M_AXI_MCU_LSU_AWID,
    output wire [              31:0] M_AXI_MCU_LSU_AWADDR,
    output wire [               3:0] M_AXI_MCU_LSU_AWREGION,
    output wire [               7:0] M_AXI_MCU_LSU_AWLEN,
    output wire [               2:0] M_AXI_MCU_LSU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_AWBURST,
    output wire                      M_AXI_MCU_LSU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_AWPROT,
    output wire [               3:0] M_AXI_MCU_LSU_AWQOS,

    output wire                      M_AXI_MCU_LSU_WVALID,
    input  wire                      M_AXI_MCU_LSU_WREADY,
    output wire [63:0]               M_AXI_MCU_LSU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_LSU_WSTRB,
    output wire                      M_AXI_MCU_LSU_WLAST,

    input  wire                      M_AXI_MCU_LSU_BVALID,
    output wire                      M_AXI_MCU_LSU_BREADY,
    input  wire [               1:0] M_AXI_MCU_LSU_BRESP,
    input  wire [18:0]               M_AXI_MCU_LSU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_LSU_ARVALID,
    input  wire                      M_AXI_MCU_LSU_ARREADY,
    output wire [18:0]               M_AXI_MCU_LSU_ARID,
    output wire [              31:0] M_AXI_MCU_LSU_ARADDR,
    output wire [               3:0] M_AXI_MCU_LSU_ARREGION,
    output wire [               7:0] M_AXI_MCU_LSU_ARLEN,
    output wire [               2:0] M_AXI_MCU_LSU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_ARBURST,
    output wire                      M_AXI_MCU_LSU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_ARPROT,
    output wire [               3:0] M_AXI_MCU_LSU_ARQOS,

    input  wire                      M_AXI_MCU_LSU_RVALID,
    output wire                      M_AXI_MCU_LSU_RREADY,
    input  wire [18:0]              M_AXI_MCU_LSU_RID,
    input  wire [              63:0] M_AXI_MCU_LSU_RDATA,
    input  wire [               1:0] M_AXI_MCU_LSU_RRESP,
    input  wire                      M_AXI_MCU_LSU_RLAST,

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_IFU_AWVALID,
    input  wire                      M_AXI_MCU_IFU_AWREADY,
    output wire [18:0]               M_AXI_MCU_IFU_AWID,
    output wire [              31:0] M_AXI_MCU_IFU_AWADDR,
    output wire [               3:0] M_AXI_MCU_IFU_AWREGION,
    output wire [               7:0] M_AXI_MCU_IFU_AWLEN,
    output wire [               2:0] M_AXI_MCU_IFU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_AWBURST,
    output wire                      M_AXI_MCU_IFU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_AWPROT,
    output wire [               3:0] M_AXI_MCU_IFU_AWQOS,

    output wire                      M_AXI_MCU_IFU_WVALID,
    input  wire                      M_AXI_MCU_IFU_WREADY,
    output wire [63:0]               M_AXI_MCU_IFU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_IFU_WSTRB,
    output wire                      M_AXI_MCU_IFU_WLAST,

    input  wire                      M_AXI_MCU_IFU_BVALID,
    output wire                      M_AXI_MCU_IFU_BREADY,
    input  wire [               1:0] M_AXI_MCU_IFU_BRESP,
    input  wire [18:0]               M_AXI_MCU_IFU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_IFU_ARVALID,
    input  wire                      M_AXI_MCU_IFU_ARREADY,
    output wire [18:0]               M_AXI_MCU_IFU_ARID,
    output wire [              31:0] M_AXI_MCU_IFU_ARADDR,
    output wire [               3:0] M_AXI_MCU_IFU_ARREGION,
    output wire [               7:0] M_AXI_MCU_IFU_ARLEN,
    output wire [               2:0] M_AXI_MCU_IFU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_ARBURST,
    output wire                      M_AXI_MCU_IFU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_ARPROT,
    output wire [               3:0] M_AXI_MCU_IFU_ARQOS,

    input  wire                      M_AXI_MCU_IFU_RVALID,
    output wire                      M_AXI_MCU_IFU_RREADY,
    input  wire [18:0]               M_AXI_MCU_IFU_RID,
    input  wire [              63:0] M_AXI_MCU_IFU_RDATA,
    input  wire [               1:0] M_AXI_MCU_IFU_RRESP,
    input  wire                      M_AXI_MCU_IFU_RLAST,


    //-------------------------- SB AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_SB_AWVALID,
    input  wire                      M_AXI_MCU_SB_AWREADY,
    output wire [18:0]               M_AXI_MCU_SB_AWID,
    output wire [              31:0] M_AXI_MCU_SB_AWADDR,
    output wire [               3:0] M_AXI_MCU_SB_AWREGION,
    output wire [               7:0] M_AXI_MCU_SB_AWLEN,
    output wire [               2:0] M_AXI_MCU_SB_AWSIZE,
    output wire [               1:0] M_AXI_MCU_SB_AWBURST,
    output wire                      M_AXI_MCU_SB_AWLOCK,
    output wire [               3:0] M_AXI_MCU_SB_AWCACHE,
    output wire [               2:0] M_AXI_MCU_SB_AWPROT,
    output wire [               3:0] M_AXI_MCU_SB_AWQOS,

    output wire                      M_AXI_MCU_SB_WVALID,
    input  wire                      M_AXI_MCU_SB_WREADY,
    output wire [63:0]               M_AXI_MCU_SB_WDATA,
    output wire [ 7:0]               M_AXI_MCU_SB_WSTRB,
    output wire                      M_AXI_MCU_SB_WLAST,

    input  wire                      M_AXI_MCU_SB_BVALID,
    output wire                      M_AXI_MCU_SB_BREADY,
    input  wire [               1:0] M_AXI_MCU_SB_BRESP,
    input  wire [18:0]               M_AXI_MCU_SB_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_SB_ARVALID,
    input  wire                      M_AXI_MCU_SB_ARREADY,
    output wire [18:0]               M_AXI_MCU_SB_ARID,
    output wire [              31:0] M_AXI_MCU_SB_ARADDR,
    output wire [               3:0] M_AXI_MCU_SB_ARREGION,
    output wire [               7:0] M_AXI_MCU_SB_ARLEN,
    output wire [               2:0] M_AXI_MCU_SB_ARSIZE,
    output wire [               1:0] M_AXI_MCU_SB_ARBURST,
    output wire                      M_AXI_MCU_SB_ARLOCK,
    output wire [               3:0] M_AXI_MCU_SB_ARCACHE,
    output wire [               2:0] M_AXI_MCU_SB_ARPROT,
    output wire [               3:0] M_AXI_MCU_SB_ARQOS,

    input  wire                      M_AXI_MCU_SB_RVALID,
    output wire                      M_AXI_MCU_SB_RREADY,
    input  wire [18:0]               M_AXI_MCU_SB_RID,
    input  wire [              63:0] M_AXI_MCU_SB_RDATA,
    input  wire [               1:0] M_AXI_MCU_SB_RRESP,
    input  wire                      M_AXI_MCU_SB_RLAST,

    // FPGA Realtime register AXI Interface
    input	wire                      S_AXI_WRAPPER_ARESETN,
    input	wire                      S_AXI_WRAPPER_AWVALID,
    output	wire                      S_AXI_WRAPPER_AWREADY,
    input	wire [31:0]               S_AXI_WRAPPER_AWADDR,
    input	wire [2:0]                S_AXI_WRAPPER_AWPROT,
    input	wire                      S_AXI_WRAPPER_WVALID,
    output	wire                      S_AXI_WRAPPER_WREADY,
    input	wire [31:0]               S_AXI_WRAPPER_WDATA,
    input	wire [3:0]                S_AXI_WRAPPER_WSTRB,
    output	wire                      S_AXI_WRAPPER_BVALID,
    input	wire                      S_AXI_WRAPPER_BREADY,
    output	wire [1:0]                S_AXI_WRAPPER_BRESP,
    input	wire                      S_AXI_WRAPPER_ARVALID,
    output	wire                      S_AXI_WRAPPER_ARREADY,
    input	wire [31:0]               S_AXI_WRAPPER_ARADDR,
    input	wire [2:0]                S_AXI_WRAPPER_ARPROT,
    output	wire                      S_AXI_WRAPPER_RVALID,
    input	wire                      S_AXI_WRAPPER_RREADY,
    output	wire [31:0]               S_AXI_WRAPPER_RDATA,
    output	wire [1:0]                S_AXI_WRAPPER_RRESP,
    
    // I3C
    input	wire                      S_AXI_I3C_AWVALID,
    output	wire                      S_AXI_I3C_AWREADY,
    input	wire [31:0]               S_AXI_I3C_AWADDR,
    input	wire [2:0]                S_AXI_I3C_AWPROT,
    input	wire                      S_AXI_I3C_WVALID,
    output	wire                      S_AXI_I3C_WREADY,
    input	wire [31:0]               S_AXI_I3C_WDATA,
    input	wire [3:0]                S_AXI_I3C_WSTRB,
    output	wire                      S_AXI_I3C_BVALID,
    input	wire                      S_AXI_I3C_BREADY,
    output	wire [1:0]                S_AXI_I3C_BRESP,
    input	wire                      S_AXI_I3C_ARVALID,
    output	wire                      S_AXI_I3C_ARREADY,
    input	wire [31:0]               S_AXI_I3C_ARADDR,
    input	wire [2:0]                S_AXI_I3C_ARPROT,
    output	wire                      S_AXI_I3C_RVALID,
    input	wire                      S_AXI_I3C_RREADY,
    output	wire [31:0]               S_AXI_I3C_RDATA,
    output	wire [1:0]                S_AXI_I3C_RRESP,
    
    input wire [1:0] S_AXI_I3C_ARBURST,
    input wire [2:0] S_AXI_I3C_ARSIZE,
    input wire [7:0] S_AXI_I3C_ARLEN,
    input wire [31:0] S_AXI_I3C_ARUSER,
    input wire [18:0] S_AXI_I3C_ARID,
    input wire S_AXI_I3C_ARLOCK,
    output wire [  18:0]           S_AXI_I3C_RID,
    output wire                   S_AXI_I3C_RLAST,
    input wire [             1:0] S_AXI_I3C_AWBURST,
    input wire [             2:0] S_AXI_I3C_AWSIZE,
    input wire [             7:0] S_AXI_I3C_AWLEN,
    input wire [31:0] S_AXI_I3C_AWUSER,
    input wire [  18:0] S_AXI_I3C_AWID,
    input wire                    S_AXI_I3C_AWLOCK,
    input  wire                  S_AXI_I3C_WLAST,
    output wire [18:0] S_AXI_I3C_BID,

// TODO: Remove
//`ifdef I3C_OUTSIDE
//    input  wire scl_i,
//    input  wire sda_i,
//    output wire scl_o,
//    output wire sda_o,
//    output wire sel_od_pp_o,
//`else
//    inout  wire i3c_scl_io,
//    inout  wire i3c_sda_io,
//`endif
    output SDA_UP,
    output SDA_PUSH,
    output SDA_PULL,
    input  SDA,
    output SCL_UP,
    output SCL_PUSH,
    output SCL_PULL,
    input  SCL,

    // SS IMEM AXI Interface
    input  wire ss_axi_bram_clk,
    input  wire ss_axi_bram_en,
    input  wire [3:0] ss_axi_bram_we,
    input  wire [15:0] ss_axi_bram_addr,
    input  wire [31:0] ss_axi_bram_din,
    output wire [31:0] ss_axi_bram_dout,
    input  wire ss_axi_bram_rst
    );

caliptra_ss_top_fpga ss_wrapper (
    
    .core_clk(core_clk),

    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_LSU_AWVALID(M_AXI_MCU_LSU_AWVALID),
    .M_AXI_MCU_LSU_AWREADY(M_AXI_MCU_LSU_AWREADY),
    .M_AXI_MCU_LSU_AWID(M_AXI_MCU_LSU_AWID),
    .M_AXI_MCU_LSU_AWADDR(M_AXI_MCU_LSU_AWADDR),
    .M_AXI_MCU_LSU_AWREGION(M_AXI_MCU_LSU_AWREGION),
    .M_AXI_MCU_LSU_AWLEN(M_AXI_MCU_LSU_AWLEN),
    .M_AXI_MCU_LSU_AWSIZE(M_AXI_MCU_LSU_AWSIZE),
    .M_AXI_MCU_LSU_AWBURST(M_AXI_MCU_LSU_AWBURST),
    .M_AXI_MCU_LSU_AWLOCK(M_AXI_MCU_LSU_AWLOCK),
    .M_AXI_MCU_LSU_AWCACHE(M_AXI_MCU_LSU_AWCACHE),
    .M_AXI_MCU_LSU_AWPROT(M_AXI_MCU_LSU_AWPROT),
    .M_AXI_MCU_LSU_AWQOS(M_AXI_MCU_LSU_AWQOS),

    .M_AXI_MCU_LSU_WVALID(M_AXI_MCU_LSU_WVALID),
    .M_AXI_MCU_LSU_WREADY(M_AXI_MCU_LSU_WREADY),
    .M_AXI_MCU_LSU_WDATA(M_AXI_MCU_LSU_WDATA),
    .M_AXI_MCU_LSU_WSTRB(M_AXI_MCU_LSU_WSTRB),
    .M_AXI_MCU_LSU_WLAST(M_AXI_MCU_LSU_WLAST),

    .M_AXI_MCU_LSU_BVALID(M_AXI_MCU_LSU_BVALID),
    .M_AXI_MCU_LSU_BREADY(M_AXI_MCU_LSU_BREADY),
    .M_AXI_MCU_LSU_BRESP(M_AXI_MCU_LSU_BRESP),
    .M_AXI_MCU_LSU_BID(M_AXI_MCU_LSU_BID),

    // AXI Read Channels
    .M_AXI_MCU_LSU_ARVALID(M_AXI_MCU_LSU_ARVALID),
    .M_AXI_MCU_LSU_ARREADY(M_AXI_MCU_LSU_ARREADY),
    .M_AXI_MCU_LSU_ARID(M_AXI_MCU_LSU_ARID),
    .M_AXI_MCU_LSU_ARADDR(M_AXI_MCU_LSU_ARADDR),
    .M_AXI_MCU_LSU_ARREGION(M_AXI_MCU_LSU_ARREGION),
    .M_AXI_MCU_LSU_ARLEN(M_AXI_MCU_LSU_ARLEN),
    .M_AXI_MCU_LSU_ARSIZE(M_AXI_MCU_LSU_ARSIZE),
    .M_AXI_MCU_LSU_ARBURST(M_AXI_MCU_LSU_ARBURST),
    .M_AXI_MCU_LSU_ARLOCK(M_AXI_MCU_LSU_ARLOCK),
    .M_AXI_MCU_LSU_ARCACHE(M_AXI_MCU_LSU_ARCACHE),
    .M_AXI_MCU_LSU_ARPROT(M_AXI_MCU_LSU_ARPROT),
    .M_AXI_MCU_LSU_ARQOS(M_AXI_MCU_LSU_ARQOS),

    .M_AXI_MCU_LSU_RVALID(M_AXI_MCU_LSU_RVALID),
    .M_AXI_MCU_LSU_RREADY(M_AXI_MCU_LSU_RREADY),
    .M_AXI_MCU_LSU_RID(M_AXI_MCU_LSU_RID),
    .M_AXI_MCU_LSU_RDATA(M_AXI_MCU_LSU_RDATA),
    .M_AXI_MCU_LSU_RRESP(M_AXI_MCU_LSU_RRESP),
    .M_AXI_MCU_LSU_RLAST(M_AXI_MCU_LSU_RLAST),

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_IFU_AWVALID(M_AXI_MCU_IFU_AWVALID),
    .M_AXI_MCU_IFU_AWREADY(M_AXI_MCU_IFU_AWREADY),
    .M_AXI_MCU_IFU_AWID(M_AXI_MCU_IFU_AWID),
    .M_AXI_MCU_IFU_AWADDR(M_AXI_MCU_IFU_AWADDR),
    .M_AXI_MCU_IFU_AWREGION(M_AXI_MCU_IFU_AWREGION),
    .M_AXI_MCU_IFU_AWLEN(M_AXI_MCU_IFU_AWLEN),
    .M_AXI_MCU_IFU_AWSIZE(M_AXI_MCU_IFU_AWSIZE),
    .M_AXI_MCU_IFU_AWBURST(M_AXI_MCU_IFU_AWBURST),
    .M_AXI_MCU_IFU_AWLOCK(M_AXI_MCU_IFU_AWLOCK),
    .M_AXI_MCU_IFU_AWCACHE(M_AXI_MCU_IFU_AWCACHE),
    .M_AXI_MCU_IFU_AWPROT(M_AXI_MCU_IFU_AWPROT),
    .M_AXI_MCU_IFU_AWQOS(M_AXI_MCU_IFU_AWQOS),

    .M_AXI_MCU_IFU_WVALID(M_AXI_MCU_IFU_WVALID),
    .M_AXI_MCU_IFU_WREADY(M_AXI_MCU_IFU_WREADY),
    .M_AXI_MCU_IFU_WDATA(M_AXI_MCU_IFU_WDATA),
    .M_AXI_MCU_IFU_WSTRB(M_AXI_MCU_IFU_WSTRB),
    .M_AXI_MCU_IFU_WLAST(M_AXI_MCU_IFU_WLAST),

    .M_AXI_MCU_IFU_BVALID(M_AXI_MCU_IFU_BVALID),
    .M_AXI_MCU_IFU_BREADY(M_AXI_MCU_IFU_BREADY),
    .M_AXI_MCU_IFU_BRESP(M_AXI_MCU_IFU_BRESP),
    .M_AXI_MCU_IFU_BID(M_AXI_MCU_IFU_BID),

    // AXI Read Channels
    .M_AXI_MCU_IFU_ARVALID(M_AXI_MCU_IFU_ARVALID),
    .M_AXI_MCU_IFU_ARREADY(M_AXI_MCU_IFU_ARREADY),
    .M_AXI_MCU_IFU_ARID(M_AXI_MCU_IFU_ARID),
    .M_AXI_MCU_IFU_ARADDR(M_AXI_MCU_IFU_ARADDR),
    .M_AXI_MCU_IFU_ARREGION(M_AXI_MCU_IFU_ARREGION),
    .M_AXI_MCU_IFU_ARLEN(M_AXI_MCU_IFU_ARLEN),
    .M_AXI_MCU_IFU_ARSIZE(M_AXI_MCU_IFU_ARSIZE),
    .M_AXI_MCU_IFU_ARBURST(M_AXI_MCU_IFU_ARBURST),
    .M_AXI_MCU_IFU_ARLOCK(M_AXI_MCU_IFU_ARLOCK),
    .M_AXI_MCU_IFU_ARCACHE(M_AXI_MCU_IFU_ARCACHE),
    .M_AXI_MCU_IFU_ARPROT(M_AXI_MCU_IFU_ARPROT),
    .M_AXI_MCU_IFU_ARQOS(M_AXI_MCU_IFU_ARQOS),

    .M_AXI_MCU_IFU_RVALID(M_AXI_MCU_IFU_RVALID),
    .M_AXI_MCU_IFU_RREADY(M_AXI_MCU_IFU_RREADY),
    .M_AXI_MCU_IFU_RID(M_AXI_MCU_IFU_RID),
    .M_AXI_MCU_IFU_RDATA(M_AXI_MCU_IFU_RDATA),
    .M_AXI_MCU_IFU_RRESP(M_AXI_MCU_IFU_RRESP),
    .M_AXI_MCU_IFU_RLAST(M_AXI_MCU_IFU_RLAST),

    //-------------------------- MCU SB AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_SB_AWVALID(M_AXI_MCU_SB_AWVALID),
    .M_AXI_MCU_SB_AWREADY(M_AXI_MCU_SB_AWREADY),
    .M_AXI_MCU_SB_AWID(M_AXI_MCU_SB_AWID),
    .M_AXI_MCU_SB_AWADDR(M_AXI_MCU_SB_AWADDR),
    .M_AXI_MCU_SB_AWREGION(M_AXI_MCU_SB_AWREGION),
    .M_AXI_MCU_SB_AWLEN(M_AXI_MCU_SB_AWLEN),
    .M_AXI_MCU_SB_AWSIZE(M_AXI_MCU_SB_AWSIZE),
    .M_AXI_MCU_SB_AWBURST(M_AXI_MCU_SB_AWBURST),
    .M_AXI_MCU_SB_AWLOCK(M_AXI_MCU_SB_AWLOCK),
    .M_AXI_MCU_SB_AWCACHE(M_AXI_MCU_SB_AWCACHE),
    .M_AXI_MCU_SB_AWPROT(M_AXI_MCU_SB_AWPROT),
    .M_AXI_MCU_SB_AWQOS(M_AXI_MCU_SB_AWQOS),

    .M_AXI_MCU_SB_WVALID(M_AXI_MCU_SB_WVALID),
    .M_AXI_MCU_SB_WREADY(M_AXI_MCU_SB_WREADY),
    .M_AXI_MCU_SB_WDATA(M_AXI_MCU_SB_WDATA),
    .M_AXI_MCU_SB_WSTRB(M_AXI_MCU_SB_WSTRB),
    .M_AXI_MCU_SB_WLAST(M_AXI_MCU_SB_WLAST),

    .M_AXI_MCU_SB_BVALID(M_AXI_MCU_SB_BVALID),
    .M_AXI_MCU_SB_BREADY(M_AXI_MCU_SB_BREADY),
    .M_AXI_MCU_SB_BRESP(M_AXI_MCU_SB_BRESP),
    .M_AXI_MCU_SB_BID(M_AXI_MCU_SB_BID),

    // AXI Read Channels
    .M_AXI_MCU_SB_ARVALID(M_AXI_MCU_SB_ARVALID),
    .M_AXI_MCU_SB_ARREADY(M_AXI_MCU_SB_ARREADY),
    .M_AXI_MCU_SB_ARID(M_AXI_MCU_SB_ARID),
    .M_AXI_MCU_SB_ARADDR(M_AXI_MCU_SB_ARADDR),
    .M_AXI_MCU_SB_ARREGION(M_AXI_MCU_SB_ARREGION),
    .M_AXI_MCU_SB_ARLEN(M_AXI_MCU_SB_ARLEN),
    .M_AXI_MCU_SB_ARSIZE(M_AXI_MCU_SB_ARSIZE),
    .M_AXI_MCU_SB_ARBURST(M_AXI_MCU_SB_ARBURST),
    .M_AXI_MCU_SB_ARLOCK(M_AXI_MCU_SB_ARLOCK),
    .M_AXI_MCU_SB_ARCACHE(M_AXI_MCU_SB_ARCACHE),
    .M_AXI_MCU_SB_ARPROT(M_AXI_MCU_SB_ARPROT),
    .M_AXI_MCU_SB_ARQOS(M_AXI_MCU_SB_ARQOS),

    .M_AXI_MCU_SB_RVALID(M_AXI_MCU_SB_RVALID),
    .M_AXI_MCU_SB_RREADY(M_AXI_MCU_SB_RREADY),
    .M_AXI_MCU_SB_RID(M_AXI_MCU_SB_RID),
    .M_AXI_MCU_SB_RDATA(M_AXI_MCU_SB_RDATA),
    .M_AXI_MCU_SB_RRESP(M_AXI_MCU_SB_RRESP),
    .M_AXI_MCU_SB_RLAST(M_AXI_MCU_SB_RLAST),
    
    // I3C
    .S_AXI_I3C_AWVALID(S_AXI_I3C_AWVALID),
    .S_AXI_I3C_AWREADY(S_AXI_I3C_AWREADY),
    .S_AXI_I3C_AWADDR(S_AXI_I3C_AWADDR),
    .S_AXI_I3C_AWPROT(S_AXI_I3C_AWPROT),
    .S_AXI_I3C_WVALID(S_AXI_I3C_WVALID),
    .S_AXI_I3C_WREADY(S_AXI_I3C_WREADY),
    .S_AXI_I3C_WDATA(S_AXI_I3C_WDATA),
    .S_AXI_I3C_WSTRB(S_AXI_I3C_WSTRB),
    .S_AXI_I3C_BVALID(S_AXI_I3C_BVALID),
    .S_AXI_I3C_BREADY(S_AXI_I3C_BREADY),
    .S_AXI_I3C_BRESP(S_AXI_I3C_BRESP),
    .S_AXI_I3C_ARVALID(S_AXI_I3C_ARVALID),
    .S_AXI_I3C_ARREADY(S_AXI_I3C_ARREADY),
    .S_AXI_I3C_ARADDR(S_AXI_I3C_ARADDR),
    .S_AXI_I3C_ARPROT(S_AXI_I3C_ARPROT),
    .S_AXI_I3C_RVALID(S_AXI_I3C_RVALID),
    .S_AXI_I3C_RREADY(S_AXI_I3C_RREADY),
    .S_AXI_I3C_RDATA(S_AXI_I3C_RDATA),
    .S_AXI_I3C_RRESP(S_AXI_I3C_RRESP),
    .S_AXI_I3C_ARBURST(S_AXI_I3C_ARBURST),
    .S_AXI_I3C_ARSIZE(S_AXI_I3C_ARSIZE),
    .S_AXI_I3C_ARLEN(S_AXI_I3C_ARLEN),
    .S_AXI_I3C_ARUSER(S_AXI_I3C_ARUSER),
    .S_AXI_I3C_ARID(S_AXI_I3C_ARID),
    .S_AXI_I3C_ARLOCK(S_AXI_I3C_ARLOCK),
    .S_AXI_I3C_RID(S_AXI_I3C_RID),
    .S_AXI_I3C_RLAST(S_AXI_I3C_RLAST),
    .S_AXI_I3C_AWBURST(S_AXI_I3C_AWBURST),
    .S_AXI_I3C_AWSIZE(S_AXI_I3C_AWSIZE),
    .S_AXI_I3C_AWLEN(S_AXI_I3C_AWLEN),
    .S_AXI_I3C_AWUSER(S_AXI_I3C_AWUSER),
    .S_AXI_I3C_AWID(S_AXI_I3C_AWID),
    .S_AXI_I3C_AWLOCK(S_AXI_I3C_AWLOCK),
    .S_AXI_I3C_WLAST(S_AXI_I3C_WLAST),
    .S_AXI_I3C_BID(S_AXI_I3C_BID),

//`ifdef I3C_OUTSIDE
//    .scl_i(scl_i),
//    .sda_i(sda_i),
//    .scl_o(scl_o),
//    .sda_o(sda_o),
//    .sel_od_pp_o(sel_od_pp_o),
//`else
//    .i3c_scl_io(i3c_scl_io),
//    .i3c_sda_io(i3c_sda_io),
//`endif

    .SDA_UP(SDA_UP),
    .SDA_PUSH(SDA_PUSH),
    .SDA_PULL(SDA_PULL),
    .SDA(SDA),
    .SCL_UP(SCL_UP),
    .SCL_PUSH(SCL_PUSH),
    .SCL_PULL(SCL_PULL),
    .SCL(SCL),

    // SS IMEM AXI Interface
    .ss_axi_bram_clk(ss_axi_bram_clk),
    .ss_axi_bram_en(ss_axi_bram_en),
    .ss_axi_bram_we(ss_axi_bram_we),
    .ss_axi_bram_addr(ss_axi_bram_addr),
    .ss_axi_bram_din(ss_axi_bram_din),
    .ss_axi_bram_dout(ss_axi_bram_dout),
    .ss_axi_bram_rst(ss_axi_bram_rst)
);

endmodule