// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef SOC_ADDRESS_MAP_DEFINES_HEADER
`define SOC_ADDRESS_MAP_DEFINES_HEADER


`define SOC_BASE_ADDR                                                                               (32'h0)
`define SOC_I3CCSR_BASE_ADDR                                                                        (32'h20004000)
`define SOC_I3CCSR_I3CBASE_START                                                                    (32'h20004000)
`define SOC_I3CCSR_I3CBASE_HCI_VERSION                                                              (32'h20004000)
`define SOC_I3CCSR_I3CBASE_HC_CONTROL                                                               (32'h20004004)
`define SOC_I3CCSR_I3CBASE_CONTROLLER_DEVICE_ADDR                                                   (32'h20004008)
`define SOC_I3CCSR_I3CBASE_HC_CAPABILITIES                                                          (32'h2000400c)
`define SOC_I3CCSR_I3CBASE_RESET_CONTROL                                                            (32'h20004010)
`define SOC_I3CCSR_I3CBASE_PRESENT_STATE                                                            (32'h20004014)
`define SOC_I3CCSR_I3CBASE_INTR_STATUS                                                              (32'h20004020)
`define SOC_I3CCSR_I3CBASE_INTR_STATUS_ENABLE                                                       (32'h20004024)
`define SOC_I3CCSR_I3CBASE_INTR_SIGNAL_ENABLE                                                       (32'h20004028)
`define SOC_I3CCSR_I3CBASE_INTR_FORCE                                                               (32'h2000402c)
`define SOC_I3CCSR_I3CBASE_DAT_SECTION_OFFSET                                                       (32'h20004030)
`define SOC_I3CCSR_I3CBASE_DCT_SECTION_OFFSET                                                       (32'h20004034)
`define SOC_I3CCSR_I3CBASE_RING_HEADERS_SECTION_OFFSET                                              (32'h20004038)
`define SOC_I3CCSR_I3CBASE_PIO_SECTION_OFFSET                                                       (32'h2000403c)
`define SOC_I3CCSR_I3CBASE_EXT_CAPS_SECTION_OFFSET                                                  (32'h20004040)
`define SOC_I3CCSR_I3CBASE_INT_CTRL_CMDS_EN                                                         (32'h2000404c)
`define SOC_I3CCSR_I3CBASE_IBI_NOTIFY_CTRL                                                          (32'h20004058)
`define SOC_I3CCSR_I3CBASE_IBI_DATA_ABORT_CTRL                                                      (32'h2000405c)
`define SOC_I3CCSR_I3CBASE_DEV_CTX_BASE_LO                                                          (32'h20004060)
`define SOC_I3CCSR_I3CBASE_DEV_CTX_BASE_HI                                                          (32'h20004064)
`define SOC_I3CCSR_I3CBASE_DEV_CTX_SG                                                               (32'h20004068)
`define SOC_I3CCSR_PIOCONTROL_START                                                                 (32'h20004080)
`define SOC_I3CCSR_PIOCONTROL_COMMAND_PORT                                                          (32'h20004080)
`define SOC_I3CCSR_PIOCONTROL_RESPONSE_PORT                                                         (32'h20004084)
`define SOC_I3CCSR_PIOCONTROL_TX_DATA_PORT                                                          (32'h20004088)
`define SOC_I3CCSR_PIOCONTROL_RX_DATA_PORT                                                          (32'h20004088)
`define SOC_I3CCSR_PIOCONTROL_IBI_PORT                                                              (32'h2000408c)
`define SOC_I3CCSR_PIOCONTROL_QUEUE_THLD_CTRL                                                       (32'h20004090)
`define SOC_I3CCSR_PIOCONTROL_DATA_BUFFER_THLD_CTRL                                                 (32'h20004094)
`define SOC_I3CCSR_PIOCONTROL_QUEUE_SIZE                                                            (32'h20004098)
`define SOC_I3CCSR_PIOCONTROL_ALT_QUEUE_SIZE                                                        (32'h2000409c)
`define SOC_I3CCSR_PIOCONTROL_PIO_INTR_STATUS                                                       (32'h200040a0)
`define SOC_I3CCSR_PIOCONTROL_PIO_INTR_STATUS_ENABLE                                                (32'h200040a4)
`define SOC_I3CCSR_PIOCONTROL_PIO_INTR_SIGNAL_ENABLE                                                (32'h200040a8)
`define SOC_I3CCSR_PIOCONTROL_PIO_INTR_FORCE                                                        (32'h200040ac)
`define SOC_I3CCSR_PIOCONTROL_PIO_CONTROL                                                           (32'h200040b0)
`define SOC_I3CCSR_I3C_EC_START                                                                     (32'h20004100)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_START                                                     (32'h20004100)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_EXTCAP_HEADER                                             (32'h20004100)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_PROT_CAP_0                                                (32'h20004104)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_PROT_CAP_1                                                (32'h20004108)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_PROT_CAP_2                                                (32'h2000410c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_PROT_CAP_3                                                (32'h20004110)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_0                                               (32'h20004114)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_1                                               (32'h20004118)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_2                                               (32'h2000411c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_3                                               (32'h20004120)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_4                                               (32'h20004124)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_5                                               (32'h20004128)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_ID_6                                               (32'h2000412c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_STATUS_0                                           (32'h20004130)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_STATUS_1                                           (32'h20004134)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_DEVICE_RESET                                              (32'h20004138)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_RECOVERY_CTRL                                             (32'h2000413c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_RECOVERY_STATUS                                           (32'h20004140)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_HW_STATUS                                                 (32'h20004144)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_CTRL_0                                      (32'h20004148)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_CTRL_1                                      (32'h2000414c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_0                                    (32'h20004150)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_1                                    (32'h20004154)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_2                                    (32'h20004158)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_3                                    (32'h2000415c)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_4                                    (32'h20004160)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_STATUS_5                                    (32'h20004164)
`define SOC_I3CCSR_I3C_EC_SECFWRECOVERYIF_INDIRECT_FIFO_DATA                                        (32'h20004168)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_START                                                       (32'h20004180)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_EXTCAP_HEADER                                               (32'h20004180)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_CONTROL                                             (32'h20004184)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_DEVICE_ADDR                                         (32'h20004188)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_CAPABILITIES                                        (32'h2000418c)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE___RSVD_0                                                    (32'h20004190)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_STATUS                                              (32'h20004194)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_DEVICE_CHAR                                         (32'h20004198)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_DEVICE_PID_LO                                       (32'h2000419c)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_INTR_STATUS                                         (32'h200041a0)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE___RSVD_1                                                    (32'h200041a4)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_INTR_SIGNAL_ENABLE                                  (32'h200041a8)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_INTR_FORCE                                          (32'h200041ac)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_CCC_CONFIG_GETCAPS                                  (32'h200041b0)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_CCC_CONFIG_RSTACT_PARAMS                            (32'h200041b4)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE_STBY_CR_VIRT_DEVICE_ADDR                                    (32'h200041b8)
`define SOC_I3CCSR_I3C_EC_STDBYCTRLMODE___RSVD_3                                                    (32'h200041bc)
`define SOC_I3CCSR_I3C_EC_TTI_START                                                                 (32'h200041c0)
`define SOC_I3CCSR_I3C_EC_TTI_EXTCAP_HEADER                                                         (32'h200041c0)
`define SOC_I3CCSR_I3C_EC_TTI_CONTROL                                                               (32'h200041c4)
`define SOC_I3CCSR_I3C_EC_TTI_STATUS                                                                (32'h200041c8)
`define SOC_I3CCSR_I3C_EC_TTI_RESET_CONTROL                                                         (32'h200041cc)
`define SOC_I3CCSR_I3C_EC_TTI_INTERRUPT_STATUS                                                      (32'h200041d0)
`define SOC_I3CCSR_I3C_EC_TTI_INTERRUPT_ENABLE                                                      (32'h200041d4)
`define SOC_I3CCSR_I3C_EC_TTI_INTERRUPT_FORCE                                                       (32'h200041d8)
`define SOC_I3CCSR_I3C_EC_TTI_RX_DESC_QUEUE_PORT                                                    (32'h200041dc)
`define SOC_I3CCSR_I3C_EC_TTI_RX_DATA_PORT                                                          (32'h200041e0)
`define SOC_I3CCSR_I3C_EC_TTI_TX_DESC_QUEUE_PORT                                                    (32'h200041e4)
`define SOC_I3CCSR_I3C_EC_TTI_TX_DATA_PORT                                                          (32'h200041e8)
`define SOC_I3CCSR_I3C_EC_TTI_IBI_PORT                                                              (32'h200041ec)
`define SOC_I3CCSR_I3C_EC_TTI_QUEUE_SIZE                                                            (32'h200041f0)
`define SOC_I3CCSR_I3C_EC_TTI_IBI_QUEUE_SIZE                                                        (32'h200041f4)
`define SOC_I3CCSR_I3C_EC_TTI_QUEUE_THLD_CTRL                                                       (32'h200041f8)
`define SOC_I3CCSR_I3C_EC_TTI_DATA_BUFFER_THLD_CTRL                                                 (32'h200041fc)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_START                                                           (32'h20004200)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_EXTCAP_HEADER                                                   (32'h20004200)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_CONTROL                                                (32'h20004204)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_STATUS                                                 (32'h20004208)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_RSVD_0                                                 (32'h2000420c)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_RSVD_1                                                 (32'h20004210)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_RSVD_2                                                 (32'h20004214)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_RSVD_3                                                 (32'h20004218)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_PAD_CONF                                                    (32'h2000421c)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_PAD_ATTR                                                    (32'h20004220)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_FEATURE_2                                              (32'h20004224)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_SOC_MGMT_FEATURE_3                                              (32'h20004228)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_R_REG                                                         (32'h2000422c)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_F_REG                                                         (32'h20004230)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_SU_DAT_REG                                                    (32'h20004234)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_HD_DAT_REG                                                    (32'h20004238)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_HIGH_REG                                                      (32'h2000423c)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_LOW_REG                                                       (32'h20004240)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_HD_STA_REG                                                    (32'h20004244)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_SU_STA_REG                                                    (32'h20004248)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_SU_STO_REG                                                    (32'h2000424c)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_FREE_REG                                                      (32'h20004250)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_AVAL_REG                                                      (32'h20004254)
`define SOC_I3CCSR_I3C_EC_SOCMGMTIF_T_IDLE_REG                                                      (32'h20004258)
`define SOC_I3CCSR_I3C_EC_CTRLCFG_START                                                             (32'h20004260)
`define SOC_I3CCSR_I3C_EC_CTRLCFG_EXTCAP_HEADER                                                     (32'h20004260)
`define SOC_I3CCSR_I3C_EC_CTRLCFG_CONTROLLER_CONFIG                                                 (32'h20004264)
`define SOC_I3CCSR_I3C_EC_TERMINATION_EXTCAP_HEADER                                                 (32'h20004268)
`define SOC_I3CCSR_DAT_BASE_ADDR                                                                    (32'h20004400)
`define SOC_I3CCSR_DAT_END_ADDR                                                                     (32'h200047ff)
`define SOC_I3CCSR_DAT_DAT_MEMORY_0                                                                 (32'h20004400)
`define SOC_I3CCSR_DAT_DAT_MEMORY_1                                                                 (32'h20004408)
`define SOC_I3CCSR_DAT_DAT_MEMORY_2                                                                 (32'h20004410)
`define SOC_I3CCSR_DAT_DAT_MEMORY_3                                                                 (32'h20004418)
`define SOC_I3CCSR_DAT_DAT_MEMORY_4                                                                 (32'h20004420)
`define SOC_I3CCSR_DAT_DAT_MEMORY_5                                                                 (32'h20004428)
`define SOC_I3CCSR_DAT_DAT_MEMORY_6                                                                 (32'h20004430)
`define SOC_I3CCSR_DAT_DAT_MEMORY_7                                                                 (32'h20004438)
`define SOC_I3CCSR_DAT_DAT_MEMORY_8                                                                 (32'h20004440)
`define SOC_I3CCSR_DAT_DAT_MEMORY_9                                                                 (32'h20004448)
`define SOC_I3CCSR_DAT_DAT_MEMORY_10                                                                (32'h20004450)
`define SOC_I3CCSR_DAT_DAT_MEMORY_11                                                                (32'h20004458)
`define SOC_I3CCSR_DAT_DAT_MEMORY_12                                                                (32'h20004460)
`define SOC_I3CCSR_DAT_DAT_MEMORY_13                                                                (32'h20004468)
`define SOC_I3CCSR_DAT_DAT_MEMORY_14                                                                (32'h20004470)
`define SOC_I3CCSR_DAT_DAT_MEMORY_15                                                                (32'h20004478)
`define SOC_I3CCSR_DAT_DAT_MEMORY_16                                                                (32'h20004480)
`define SOC_I3CCSR_DAT_DAT_MEMORY_17                                                                (32'h20004488)
`define SOC_I3CCSR_DAT_DAT_MEMORY_18                                                                (32'h20004490)
`define SOC_I3CCSR_DAT_DAT_MEMORY_19                                                                (32'h20004498)
`define SOC_I3CCSR_DAT_DAT_MEMORY_20                                                                (32'h200044a0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_21                                                                (32'h200044a8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_22                                                                (32'h200044b0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_23                                                                (32'h200044b8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_24                                                                (32'h200044c0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_25                                                                (32'h200044c8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_26                                                                (32'h200044d0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_27                                                                (32'h200044d8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_28                                                                (32'h200044e0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_29                                                                (32'h200044e8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_30                                                                (32'h200044f0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_31                                                                (32'h200044f8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_32                                                                (32'h20004500)
`define SOC_I3CCSR_DAT_DAT_MEMORY_33                                                                (32'h20004508)
`define SOC_I3CCSR_DAT_DAT_MEMORY_34                                                                (32'h20004510)
`define SOC_I3CCSR_DAT_DAT_MEMORY_35                                                                (32'h20004518)
`define SOC_I3CCSR_DAT_DAT_MEMORY_36                                                                (32'h20004520)
`define SOC_I3CCSR_DAT_DAT_MEMORY_37                                                                (32'h20004528)
`define SOC_I3CCSR_DAT_DAT_MEMORY_38                                                                (32'h20004530)
`define SOC_I3CCSR_DAT_DAT_MEMORY_39                                                                (32'h20004538)
`define SOC_I3CCSR_DAT_DAT_MEMORY_40                                                                (32'h20004540)
`define SOC_I3CCSR_DAT_DAT_MEMORY_41                                                                (32'h20004548)
`define SOC_I3CCSR_DAT_DAT_MEMORY_42                                                                (32'h20004550)
`define SOC_I3CCSR_DAT_DAT_MEMORY_43                                                                (32'h20004558)
`define SOC_I3CCSR_DAT_DAT_MEMORY_44                                                                (32'h20004560)
`define SOC_I3CCSR_DAT_DAT_MEMORY_45                                                                (32'h20004568)
`define SOC_I3CCSR_DAT_DAT_MEMORY_46                                                                (32'h20004570)
`define SOC_I3CCSR_DAT_DAT_MEMORY_47                                                                (32'h20004578)
`define SOC_I3CCSR_DAT_DAT_MEMORY_48                                                                (32'h20004580)
`define SOC_I3CCSR_DAT_DAT_MEMORY_49                                                                (32'h20004588)
`define SOC_I3CCSR_DAT_DAT_MEMORY_50                                                                (32'h20004590)
`define SOC_I3CCSR_DAT_DAT_MEMORY_51                                                                (32'h20004598)
`define SOC_I3CCSR_DAT_DAT_MEMORY_52                                                                (32'h200045a0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_53                                                                (32'h200045a8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_54                                                                (32'h200045b0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_55                                                                (32'h200045b8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_56                                                                (32'h200045c0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_57                                                                (32'h200045c8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_58                                                                (32'h200045d0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_59                                                                (32'h200045d8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_60                                                                (32'h200045e0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_61                                                                (32'h200045e8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_62                                                                (32'h200045f0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_63                                                                (32'h200045f8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_64                                                                (32'h20004600)
`define SOC_I3CCSR_DAT_DAT_MEMORY_65                                                                (32'h20004608)
`define SOC_I3CCSR_DAT_DAT_MEMORY_66                                                                (32'h20004610)
`define SOC_I3CCSR_DAT_DAT_MEMORY_67                                                                (32'h20004618)
`define SOC_I3CCSR_DAT_DAT_MEMORY_68                                                                (32'h20004620)
`define SOC_I3CCSR_DAT_DAT_MEMORY_69                                                                (32'h20004628)
`define SOC_I3CCSR_DAT_DAT_MEMORY_70                                                                (32'h20004630)
`define SOC_I3CCSR_DAT_DAT_MEMORY_71                                                                (32'h20004638)
`define SOC_I3CCSR_DAT_DAT_MEMORY_72                                                                (32'h20004640)
`define SOC_I3CCSR_DAT_DAT_MEMORY_73                                                                (32'h20004648)
`define SOC_I3CCSR_DAT_DAT_MEMORY_74                                                                (32'h20004650)
`define SOC_I3CCSR_DAT_DAT_MEMORY_75                                                                (32'h20004658)
`define SOC_I3CCSR_DAT_DAT_MEMORY_76                                                                (32'h20004660)
`define SOC_I3CCSR_DAT_DAT_MEMORY_77                                                                (32'h20004668)
`define SOC_I3CCSR_DAT_DAT_MEMORY_78                                                                (32'h20004670)
`define SOC_I3CCSR_DAT_DAT_MEMORY_79                                                                (32'h20004678)
`define SOC_I3CCSR_DAT_DAT_MEMORY_80                                                                (32'h20004680)
`define SOC_I3CCSR_DAT_DAT_MEMORY_81                                                                (32'h20004688)
`define SOC_I3CCSR_DAT_DAT_MEMORY_82                                                                (32'h20004690)
`define SOC_I3CCSR_DAT_DAT_MEMORY_83                                                                (32'h20004698)
`define SOC_I3CCSR_DAT_DAT_MEMORY_84                                                                (32'h200046a0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_85                                                                (32'h200046a8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_86                                                                (32'h200046b0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_87                                                                (32'h200046b8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_88                                                                (32'h200046c0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_89                                                                (32'h200046c8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_90                                                                (32'h200046d0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_91                                                                (32'h200046d8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_92                                                                (32'h200046e0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_93                                                                (32'h200046e8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_94                                                                (32'h200046f0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_95                                                                (32'h200046f8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_96                                                                (32'h20004700)
`define SOC_I3CCSR_DAT_DAT_MEMORY_97                                                                (32'h20004708)
`define SOC_I3CCSR_DAT_DAT_MEMORY_98                                                                (32'h20004710)
`define SOC_I3CCSR_DAT_DAT_MEMORY_99                                                                (32'h20004718)
`define SOC_I3CCSR_DAT_DAT_MEMORY_100                                                               (32'h20004720)
`define SOC_I3CCSR_DAT_DAT_MEMORY_101                                                               (32'h20004728)
`define SOC_I3CCSR_DAT_DAT_MEMORY_102                                                               (32'h20004730)
`define SOC_I3CCSR_DAT_DAT_MEMORY_103                                                               (32'h20004738)
`define SOC_I3CCSR_DAT_DAT_MEMORY_104                                                               (32'h20004740)
`define SOC_I3CCSR_DAT_DAT_MEMORY_105                                                               (32'h20004748)
`define SOC_I3CCSR_DAT_DAT_MEMORY_106                                                               (32'h20004750)
`define SOC_I3CCSR_DAT_DAT_MEMORY_107                                                               (32'h20004758)
`define SOC_I3CCSR_DAT_DAT_MEMORY_108                                                               (32'h20004760)
`define SOC_I3CCSR_DAT_DAT_MEMORY_109                                                               (32'h20004768)
`define SOC_I3CCSR_DAT_DAT_MEMORY_110                                                               (32'h20004770)
`define SOC_I3CCSR_DAT_DAT_MEMORY_111                                                               (32'h20004778)
`define SOC_I3CCSR_DAT_DAT_MEMORY_112                                                               (32'h20004780)
`define SOC_I3CCSR_DAT_DAT_MEMORY_113                                                               (32'h20004788)
`define SOC_I3CCSR_DAT_DAT_MEMORY_114                                                               (32'h20004790)
`define SOC_I3CCSR_DAT_DAT_MEMORY_115                                                               (32'h20004798)
`define SOC_I3CCSR_DAT_DAT_MEMORY_116                                                               (32'h200047a0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_117                                                               (32'h200047a8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_118                                                               (32'h200047b0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_119                                                               (32'h200047b8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_120                                                               (32'h200047c0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_121                                                               (32'h200047c8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_122                                                               (32'h200047d0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_123                                                               (32'h200047d8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_124                                                               (32'h200047e0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_125                                                               (32'h200047e8)
`define SOC_I3CCSR_DAT_DAT_MEMORY_126                                                               (32'h200047f0)
`define SOC_I3CCSR_DAT_DAT_MEMORY_127                                                               (32'h200047f8)
`define SOC_I3CCSR_DCT_BASE_ADDR                                                                    (32'h20004800)
`define SOC_I3CCSR_DCT_END_ADDR                                                                     (32'h20004fff)
`define SOC_I3CCSR_DCT_DCT_MEMORY_0                                                                 (32'h20004800)
`define SOC_I3CCSR_DCT_DCT_MEMORY_1                                                                 (32'h20004810)
`define SOC_I3CCSR_DCT_DCT_MEMORY_2                                                                 (32'h20004820)
`define SOC_I3CCSR_DCT_DCT_MEMORY_3                                                                 (32'h20004830)
`define SOC_I3CCSR_DCT_DCT_MEMORY_4                                                                 (32'h20004840)
`define SOC_I3CCSR_DCT_DCT_MEMORY_5                                                                 (32'h20004850)
`define SOC_I3CCSR_DCT_DCT_MEMORY_6                                                                 (32'h20004860)
`define SOC_I3CCSR_DCT_DCT_MEMORY_7                                                                 (32'h20004870)
`define SOC_I3CCSR_DCT_DCT_MEMORY_8                                                                 (32'h20004880)
`define SOC_I3CCSR_DCT_DCT_MEMORY_9                                                                 (32'h20004890)
`define SOC_I3CCSR_DCT_DCT_MEMORY_10                                                                (32'h200048a0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_11                                                                (32'h200048b0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_12                                                                (32'h200048c0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_13                                                                (32'h200048d0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_14                                                                (32'h200048e0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_15                                                                (32'h200048f0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_16                                                                (32'h20004900)
`define SOC_I3CCSR_DCT_DCT_MEMORY_17                                                                (32'h20004910)
`define SOC_I3CCSR_DCT_DCT_MEMORY_18                                                                (32'h20004920)
`define SOC_I3CCSR_DCT_DCT_MEMORY_19                                                                (32'h20004930)
`define SOC_I3CCSR_DCT_DCT_MEMORY_20                                                                (32'h20004940)
`define SOC_I3CCSR_DCT_DCT_MEMORY_21                                                                (32'h20004950)
`define SOC_I3CCSR_DCT_DCT_MEMORY_22                                                                (32'h20004960)
`define SOC_I3CCSR_DCT_DCT_MEMORY_23                                                                (32'h20004970)
`define SOC_I3CCSR_DCT_DCT_MEMORY_24                                                                (32'h20004980)
`define SOC_I3CCSR_DCT_DCT_MEMORY_25                                                                (32'h20004990)
`define SOC_I3CCSR_DCT_DCT_MEMORY_26                                                                (32'h200049a0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_27                                                                (32'h200049b0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_28                                                                (32'h200049c0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_29                                                                (32'h200049d0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_30                                                                (32'h200049e0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_31                                                                (32'h200049f0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_32                                                                (32'h20004a00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_33                                                                (32'h20004a10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_34                                                                (32'h20004a20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_35                                                                (32'h20004a30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_36                                                                (32'h20004a40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_37                                                                (32'h20004a50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_38                                                                (32'h20004a60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_39                                                                (32'h20004a70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_40                                                                (32'h20004a80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_41                                                                (32'h20004a90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_42                                                                (32'h20004aa0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_43                                                                (32'h20004ab0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_44                                                                (32'h20004ac0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_45                                                                (32'h20004ad0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_46                                                                (32'h20004ae0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_47                                                                (32'h20004af0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_48                                                                (32'h20004b00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_49                                                                (32'h20004b10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_50                                                                (32'h20004b20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_51                                                                (32'h20004b30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_52                                                                (32'h20004b40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_53                                                                (32'h20004b50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_54                                                                (32'h20004b60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_55                                                                (32'h20004b70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_56                                                                (32'h20004b80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_57                                                                (32'h20004b90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_58                                                                (32'h20004ba0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_59                                                                (32'h20004bb0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_60                                                                (32'h20004bc0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_61                                                                (32'h20004bd0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_62                                                                (32'h20004be0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_63                                                                (32'h20004bf0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_64                                                                (32'h20004c00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_65                                                                (32'h20004c10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_66                                                                (32'h20004c20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_67                                                                (32'h20004c30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_68                                                                (32'h20004c40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_69                                                                (32'h20004c50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_70                                                                (32'h20004c60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_71                                                                (32'h20004c70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_72                                                                (32'h20004c80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_73                                                                (32'h20004c90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_74                                                                (32'h20004ca0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_75                                                                (32'h20004cb0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_76                                                                (32'h20004cc0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_77                                                                (32'h20004cd0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_78                                                                (32'h20004ce0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_79                                                                (32'h20004cf0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_80                                                                (32'h20004d00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_81                                                                (32'h20004d10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_82                                                                (32'h20004d20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_83                                                                (32'h20004d30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_84                                                                (32'h20004d40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_85                                                                (32'h20004d50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_86                                                                (32'h20004d60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_87                                                                (32'h20004d70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_88                                                                (32'h20004d80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_89                                                                (32'h20004d90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_90                                                                (32'h20004da0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_91                                                                (32'h20004db0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_92                                                                (32'h20004dc0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_93                                                                (32'h20004dd0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_94                                                                (32'h20004de0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_95                                                                (32'h20004df0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_96                                                                (32'h20004e00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_97                                                                (32'h20004e10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_98                                                                (32'h20004e20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_99                                                                (32'h20004e30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_100                                                               (32'h20004e40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_101                                                               (32'h20004e50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_102                                                               (32'h20004e60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_103                                                               (32'h20004e70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_104                                                               (32'h20004e80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_105                                                               (32'h20004e90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_106                                                               (32'h20004ea0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_107                                                               (32'h20004eb0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_108                                                               (32'h20004ec0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_109                                                               (32'h20004ed0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_110                                                               (32'h20004ee0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_111                                                               (32'h20004ef0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_112                                                               (32'h20004f00)
`define SOC_I3CCSR_DCT_DCT_MEMORY_113                                                               (32'h20004f10)
`define SOC_I3CCSR_DCT_DCT_MEMORY_114                                                               (32'h20004f20)
`define SOC_I3CCSR_DCT_DCT_MEMORY_115                                                               (32'h20004f30)
`define SOC_I3CCSR_DCT_DCT_MEMORY_116                                                               (32'h20004f40)
`define SOC_I3CCSR_DCT_DCT_MEMORY_117                                                               (32'h20004f50)
`define SOC_I3CCSR_DCT_DCT_MEMORY_118                                                               (32'h20004f60)
`define SOC_I3CCSR_DCT_DCT_MEMORY_119                                                               (32'h20004f70)
`define SOC_I3CCSR_DCT_DCT_MEMORY_120                                                               (32'h20004f80)
`define SOC_I3CCSR_DCT_DCT_MEMORY_121                                                               (32'h20004f90)
`define SOC_I3CCSR_DCT_DCT_MEMORY_122                                                               (32'h20004fa0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_123                                                               (32'h20004fb0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_124                                                               (32'h20004fc0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_125                                                               (32'h20004fd0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_126                                                               (32'h20004fe0)
`define SOC_I3CCSR_DCT_DCT_MEMORY_127                                                               (32'h20004ff0)
`define SOC_MCI_REG_BASE_ADDR                                                                       (32'h21000000)
`define SOC_MCI_REG_HW_CAPABILITIES                                                                 (32'h21000000)
`define SOC_MCI_REG_FW_CAPABILITIES                                                                 (32'h21000004)
`define SOC_MCI_REG_CAP_LOCK                                                                        (32'h21000008)
`define SOC_MCI_REG_HW_REV_ID                                                                       (32'h2100000c)
`define SOC_MCI_REG_FW_REV_ID_0                                                                     (32'h21000010)
`define SOC_MCI_REG_FW_REV_ID_1                                                                     (32'h21000014)
`define SOC_MCI_REG_HW_CONFIG0                                                                      (32'h21000018)
`define SOC_MCI_REG_HW_CONFIG1                                                                      (32'h2100001c)
`define SOC_MCI_REG_FW_FLOW_STATUS                                                                  (32'h21000020)
`define SOC_MCI_REG_HW_FLOW_STATUS                                                                  (32'h21000024)
`define SOC_MCI_REG_RESET_REASON                                                                    (32'h21000028)
`define SOC_MCI_REG_RESET_STATUS                                                                    (32'h2100002c)
`define SOC_MCI_REG_SECURITY_STATE                                                                  (32'h21000030)
`define SOC_MCI_REG_HW_ERROR_FATAL                                                                  (32'h21000040)
`define SOC_MCI_REG_AGG_ERROR_FATAL                                                                 (32'h21000044)
`define SOC_MCI_REG_HW_ERROR_NON_FATAL                                                              (32'h21000048)
`define SOC_MCI_REG_AGG_ERROR_NON_FATAL                                                             (32'h2100004c)
`define SOC_MCI_REG_FW_ERROR_FATAL                                                                  (32'h21000050)
`define SOC_MCI_REG_FW_ERROR_NON_FATAL                                                              (32'h21000054)
`define SOC_MCI_REG_HW_ERROR_ENC                                                                    (32'h21000058)
`define SOC_MCI_REG_FW_ERROR_ENC                                                                    (32'h2100005c)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_0                                                        (32'h21000060)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_1                                                        (32'h21000064)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_2                                                        (32'h21000068)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_3                                                        (32'h2100006c)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_4                                                        (32'h21000070)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_5                                                        (32'h21000074)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_6                                                        (32'h21000078)
`define SOC_MCI_REG_FW_EXTENDED_ERROR_INFO_7                                                        (32'h2100007c)
`define SOC_MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                    (32'h21000080)
`define SOC_MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                                (32'h21000084)
`define SOC_MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK                                                   (32'h21000088)
`define SOC_MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK                                               (32'h2100008c)
`define SOC_MCI_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                    (32'h21000090)
`define SOC_MCI_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                                (32'h21000094)
`define SOC_MCI_REG_WDT_TIMER1_EN                                                                   (32'h210000a0)
`define SOC_MCI_REG_WDT_TIMER1_CTRL                                                                 (32'h210000a4)
`define SOC_MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_0                                                     (32'h210000a8)
`define SOC_MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_1                                                     (32'h210000ac)
`define SOC_MCI_REG_WDT_TIMER2_EN                                                                   (32'h210000b0)
`define SOC_MCI_REG_WDT_TIMER2_CTRL                                                                 (32'h210000b4)
`define SOC_MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_0                                                     (32'h210000b8)
`define SOC_MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_1                                                     (32'h210000bc)
`define SOC_MCI_REG_WDT_STATUS                                                                      (32'h210000c0)
`define SOC_MCI_REG_WDT_CFG_0                                                                       (32'h210000d0)
`define SOC_MCI_REG_WDT_CFG_1                                                                       (32'h210000d4)
`define SOC_MCI_REG_MCU_TIMER_CONFIG                                                                (32'h210000e0)
`define SOC_MCI_REG_MCU_RV_MTIME_L                                                                  (32'h210000e4)
`define SOC_MCI_REG_MCU_RV_MTIME_H                                                                  (32'h210000e8)
`define SOC_MCI_REG_MCU_RV_MTIMECMP_L                                                               (32'h210000ec)
`define SOC_MCI_REG_MCU_RV_MTIMECMP_H                                                               (32'h210000f0)
`define SOC_MCI_REG_RESET_REQUEST                                                                   (32'h21000100)
`define SOC_MCI_REG_MCI_BOOTFSM_GO                                                                  (32'h21000104)
`define SOC_MCI_REG_FW_SRAM_EXEC_REGION_SIZE                                                        (32'h21000108)
`define SOC_MCI_REG_MCU_NMI_VECTOR                                                                  (32'h2100010c)
`define SOC_MCI_REG_MCU_RESET_VECTOR                                                                (32'h21000110)
`define SOC_MCI_REG_MBOX0_VALID_AXI_USER_0                                                          (32'h21000180)
`define SOC_MCI_REG_MBOX0_VALID_AXI_USER_1                                                          (32'h21000184)
`define SOC_MCI_REG_MBOX0_VALID_AXI_USER_2                                                          (32'h21000188)
`define SOC_MCI_REG_MBOX0_VALID_AXI_USER_3                                                          (32'h2100018c)
`define SOC_MCI_REG_MBOX0_VALID_AXI_USER_4                                                          (32'h21000190)
`define SOC_MCI_REG_MBOX0_AXI_USER_LOCK_0                                                           (32'h210001a0)
`define SOC_MCI_REG_MBOX0_AXI_USER_LOCK_1                                                           (32'h210001a4)
`define SOC_MCI_REG_MBOX0_AXI_USER_LOCK_2                                                           (32'h210001a8)
`define SOC_MCI_REG_MBOX0_AXI_USER_LOCK_3                                                           (32'h210001ac)
`define SOC_MCI_REG_MBOX0_AXI_USER_LOCK_4                                                           (32'h210001b0)
`define SOC_MCI_REG_MBOX1_VALID_AXI_USER_0                                                          (32'h210001c0)
`define SOC_MCI_REG_MBOX1_VALID_AXI_USER_1                                                          (32'h210001c4)
`define SOC_MCI_REG_MBOX1_VALID_AXI_USER_2                                                          (32'h210001c8)
`define SOC_MCI_REG_MBOX1_VALID_AXI_USER_3                                                          (32'h210001cc)
`define SOC_MCI_REG_MBOX1_VALID_AXI_USER_4                                                          (32'h210001d0)
`define SOC_MCI_REG_MBOX1_AXI_USER_LOCK_0                                                           (32'h210001e0)
`define SOC_MCI_REG_MBOX1_AXI_USER_LOCK_1                                                           (32'h210001e4)
`define SOC_MCI_REG_MBOX1_AXI_USER_LOCK_2                                                           (32'h210001e8)
`define SOC_MCI_REG_MBOX1_AXI_USER_LOCK_3                                                           (32'h210001ec)
`define SOC_MCI_REG_MBOX1_AXI_USER_LOCK_4                                                           (32'h210001f0)
`define SOC_MCI_REG_GENERIC_INPUT_WIRES_0                                                           (32'h21000400)
`define SOC_MCI_REG_GENERIC_INPUT_WIRES_1                                                           (32'h21000404)
`define SOC_MCI_REG_GENERIC_OUTPUT_WIRES_0                                                          (32'h21000408)
`define SOC_MCI_REG_GENERIC_OUTPUT_WIRES_1                                                          (32'h2100040c)
`define SOC_MCI_REG_DEBUG_IN                                                                        (32'h21000410)
`define SOC_MCI_REG_DEBUG_OUT                                                                       (32'h21000414)
`define SOC_MCI_REG_SS_DEBUG_INTENT                                                                 (32'h21000418)
`define SOC_MCI_REG_SS_CONFIG_DONE                                                                  (32'h21000440)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_0                                               (32'h21000480)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_1                                               (32'h21000484)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_2                                               (32'h21000488)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_3                                               (32'h2100048c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_4                                               (32'h21000490)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_5                                               (32'h21000494)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_6                                               (32'h21000498)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_7                                               (32'h2100049c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_8                                               (32'h210004a0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_9                                               (32'h210004a4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_10                                              (32'h210004a8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_11                                              (32'h210004ac)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_0                                               (32'h210004b0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_1                                               (32'h210004b4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_2                                               (32'h210004b8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_3                                               (32'h210004bc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_4                                               (32'h210004c0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_5                                               (32'h210004c4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_6                                               (32'h210004c8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_7                                               (32'h210004cc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_8                                               (32'h210004d0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_9                                               (32'h210004d4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_10                                              (32'h210004d8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_11                                              (32'h210004dc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_0                                               (32'h210004e0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_1                                               (32'h210004e4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_2                                               (32'h210004e8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_3                                               (32'h210004ec)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_4                                               (32'h210004f0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_5                                               (32'h210004f4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_6                                               (32'h210004f8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_7                                               (32'h210004fc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_8                                               (32'h21000500)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_9                                               (32'h21000504)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_10                                              (32'h21000508)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_11                                              (32'h2100050c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_0                                               (32'h21000510)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_1                                               (32'h21000514)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_2                                               (32'h21000518)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_3                                               (32'h2100051c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_4                                               (32'h21000520)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_5                                               (32'h21000524)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_6                                               (32'h21000528)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_7                                               (32'h2100052c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_8                                               (32'h21000530)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_9                                               (32'h21000534)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_10                                              (32'h21000538)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_11                                              (32'h2100053c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_0                                               (32'h21000540)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_1                                               (32'h21000544)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_2                                               (32'h21000548)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_3                                               (32'h2100054c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_4                                               (32'h21000550)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_5                                               (32'h21000554)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_6                                               (32'h21000558)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_7                                               (32'h2100055c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_8                                               (32'h21000560)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_9                                               (32'h21000564)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_10                                              (32'h21000568)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_11                                              (32'h2100056c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_0                                               (32'h21000570)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_1                                               (32'h21000574)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_2                                               (32'h21000578)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_3                                               (32'h2100057c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_4                                               (32'h21000580)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_5                                               (32'h21000584)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_6                                               (32'h21000588)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_7                                               (32'h2100058c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_8                                               (32'h21000590)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_9                                               (32'h21000594)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_10                                              (32'h21000598)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_11                                              (32'h2100059c)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_0                                               (32'h210005a0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_1                                               (32'h210005a4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_2                                               (32'h210005a8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_3                                               (32'h210005ac)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_4                                               (32'h210005b0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_5                                               (32'h210005b4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_6                                               (32'h210005b8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_7                                               (32'h210005bc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_8                                               (32'h210005c0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_9                                               (32'h210005c4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_10                                              (32'h210005c8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_11                                              (32'h210005cc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_0                                               (32'h210005d0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_1                                               (32'h210005d4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_2                                               (32'h210005d8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_3                                               (32'h210005dc)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_4                                               (32'h210005e0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_5                                               (32'h210005e4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_6                                               (32'h210005e8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_7                                               (32'h210005ec)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_8                                               (32'h210005f0)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_9                                               (32'h210005f4)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_10                                              (32'h210005f8)
`define SOC_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_11                                              (32'h210005fc)
`define SOC_MCI_REG_INTR_BLOCK_RF_START                                                             (32'h21001000)
`define SOC_MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h21001000)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R                                                  (32'h21001004)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R                                                  (32'h21001008)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R                                                  (32'h2100100c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R                                                  (32'h21001010)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h21001014)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h21001018)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R                                            (32'h2100101c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R                                            (32'h21001020)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R                                            (32'h21001024)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R                                            (32'h21001028)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R                                                (32'h2100102c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R                                                (32'h21001030)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R                                                (32'h21001034)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R                                                (32'h21001038)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h21001100)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_INV_DEV_INTR_COUNT_R                                  (32'h21001104)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_INV_DEV_INTR_COUNT_R                                  (32'h21001108)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_CMD_FAIL_INTR_COUNT_R                                 (32'h2100110c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_CMD_FAIL_INTR_COUNT_R                                 (32'h21001110)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_ECC_UNC_INTR_COUNT_R                                  (32'h21001114)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_ECC_UNC_INTR_COUNT_R                                  (32'h21001118)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MCU_SRAM_DMI_AXI_COLLISION_INTR_COUNT_R                     (32'h2100111c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                             (32'h21001120)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                             (32'h21001124)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_R                               (32'h21001128)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_R                               (32'h2100112c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_R                               (32'h21001130)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_R                               (32'h21001134)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_R                               (32'h21001138)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_R                               (32'h2100113c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_R                               (32'h21001140)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_R                               (32'h21001144)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_R                               (32'h21001148)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_R                               (32'h2100114c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_R                              (32'h21001150)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_R                              (32'h21001154)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_R                              (32'h21001158)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_R                              (32'h2100115c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_R                              (32'h21001160)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_R                              (32'h21001164)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_R                              (32'h21001168)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_R                              (32'h2100116c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_R                              (32'h21001170)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_R                              (32'h21001174)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_R                              (32'h21001178)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_R                              (32'h2100117c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_R                              (32'h21001180)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_R                              (32'h21001184)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_R                              (32'h21001188)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_R                              (32'h2100118c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_R                              (32'h21001190)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_R                              (32'h21001194)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_R                              (32'h21001198)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_R                              (32'h2100119c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_R                              (32'h210011a0)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_R                              (32'h210011a4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_R                               (32'h21001200)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MCU_RESET_REQ_INTR_COUNT_R                            (32'h21001204)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_R                                  (32'h21001208)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_R                           (32'h2100120c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_R                           (32'h21001210)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_R                           (32'h21001214)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_R                           (32'h21001218)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_R                           (32'h2100121c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_R                           (32'h21001220)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_R                           (32'h21001224)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_R                           (32'h21001228)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_R                           (32'h2100122c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_R                           (32'h21001230)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_R                          (32'h21001234)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_R                          (32'h21001238)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_R                          (32'h2100123c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_R                          (32'h21001240)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_R                          (32'h21001244)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_R                          (32'h21001248)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_R                          (32'h2100124c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_R                          (32'h21001250)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_R                          (32'h21001254)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_R                          (32'h21001258)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_R                          (32'h2100125c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_R                          (32'h21001260)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_R                          (32'h21001264)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_R                          (32'h21001268)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_R                          (32'h2100126c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_R                          (32'h21001270)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_R                          (32'h21001274)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_R                          (32'h21001278)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_R                          (32'h2100127c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_R                          (32'h21001280)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_R                          (32'h21001284)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_R                          (32'h21001288)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_CMD_AVAIL_INTR_COUNT_R                                (32'h2100128c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_CMD_AVAIL_INTR_COUNT_R                                (32'h21001290)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_ECC_COR_INTR_COUNT_R                                  (32'h21001294)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_ECC_COR_INTR_COUNT_R                                  (32'h21001298)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                                   (32'h2100129c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_R                                      (32'h210012a0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_SOC_REQ_LOCK_INTR_COUNT_R                             (32'h210012a4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_SOC_REQ_LOCK_INTR_COUNT_R                             (32'h210012a8)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h21001300)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_INV_DEV_INTR_COUNT_INCR_R                             (32'h21001304)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_INV_DEV_INTR_COUNT_INCR_R                             (32'h21001308)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_CMD_FAIL_INTR_COUNT_INCR_R                            (32'h2100130c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_CMD_FAIL_INTR_COUNT_INCR_R                            (32'h21001310)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_ECC_UNC_INTR_COUNT_INCR_R                             (32'h21001314)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_ECC_UNC_INTR_COUNT_INCR_R                             (32'h21001318)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                        (32'h2100131c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                        (32'h21001320)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_MCU_SRAM_DMI_AXI_COLLISION_INTR_COUNT_INCR_R                (32'h21001324)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R                          (32'h21001328)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R                          (32'h2100132c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R                          (32'h21001330)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R                          (32'h21001334)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R                          (32'h21001338)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R                          (32'h2100133c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R                          (32'h21001340)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R                          (32'h21001344)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R                          (32'h21001348)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R                          (32'h2100134c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R                         (32'h21001350)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R                         (32'h21001354)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R                         (32'h21001358)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R                         (32'h2100135c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R                         (32'h21001360)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R                         (32'h21001364)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R                         (32'h21001368)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R                         (32'h2100136c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R                         (32'h21001370)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R                         (32'h21001374)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R                         (32'h21001378)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R                         (32'h2100137c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R                         (32'h21001380)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R                         (32'h21001384)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R                         (32'h21001388)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R                         (32'h2100138c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R                         (32'h21001390)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R                         (32'h21001394)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R                         (32'h21001398)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R                         (32'h2100139c)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R                         (32'h210013a0)
`define SOC_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R                         (32'h210013a4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R                          (32'h210013a8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MCU_RESET_REQ_INTR_COUNT_INCR_R                       (32'h210013ac)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R                             (32'h210013b0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R                      (32'h210013b4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R                      (32'h210013b8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R                      (32'h210013bc)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R                      (32'h210013c0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R                      (32'h210013c4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R                      (32'h210013c8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R                      (32'h210013cc)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R                      (32'h210013d0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R                      (32'h210013d4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R                      (32'h210013d8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R                     (32'h210013dc)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R                     (32'h210013e0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R                     (32'h210013e4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R                     (32'h210013e8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R                     (32'h210013ec)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R                     (32'h210013f0)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R                     (32'h210013f4)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R                     (32'h210013f8)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R                     (32'h210013fc)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R                     (32'h21001400)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R                     (32'h21001404)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R                     (32'h21001408)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R                     (32'h2100140c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R                     (32'h21001410)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R                     (32'h21001414)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R                     (32'h21001418)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R                     (32'h2100141c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R                     (32'h21001420)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R                     (32'h21001424)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R                     (32'h21001428)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R                     (32'h2100142c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R                     (32'h21001430)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_CMD_AVAIL_INTR_COUNT_INCR_R                           (32'h21001434)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_CMD_AVAIL_INTR_COUNT_INCR_R                           (32'h21001438)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_ECC_COR_INTR_COUNT_INCR_R                             (32'h2100143c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_ECC_COR_INTR_COUNT_INCR_R                             (32'h21001440)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                              (32'h21001444)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R                                 (32'h21001448)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_SOC_REQ_LOCK_INTR_COUNT_INCR_R                        (32'h2100144c)
`define SOC_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_SOC_REQ_LOCK_INTR_COUNT_INCR_R                        (32'h21001450)
`define SOC_MBOX_CSR_BASE_ADDR                                                                      (32'h30020000)
`define SOC_MBOX_CSR_MBOX_LOCK                                                                      (32'h30020000)
`define SOC_MBOX_CSR_MBOX_USER                                                                      (32'h30020004)
`define SOC_MBOX_CSR_MBOX_CMD                                                                       (32'h30020008)
`define SOC_MBOX_CSR_MBOX_DLEN                                                                      (32'h3002000c)
`define SOC_MBOX_CSR_MBOX_DATAIN                                                                    (32'h30020010)
`define SOC_MBOX_CSR_MBOX_DATAOUT                                                                   (32'h30020014)
`define SOC_MBOX_CSR_MBOX_EXECUTE                                                                   (32'h30020018)
`define SOC_MBOX_CSR_MBOX_STATUS                                                                    (32'h3002001c)
`define SOC_MBOX_CSR_MBOX_UNLOCK                                                                    (32'h30020020)
`define SOC_MBOX_CSR_TAP_MODE                                                                       (32'h30020024)
`define SOC_SHA512_ACC_CSR_BASE_ADDR                                                                (32'h30021000)
`define SOC_SHA512_ACC_CSR_LOCK                                                                     (32'h30021000)
`define SOC_SHA512_ACC_CSR_USER                                                                     (32'h30021004)
`define SOC_SHA512_ACC_CSR_MODE                                                                     (32'h30021008)
`define SOC_SHA512_ACC_CSR_START_ADDRESS                                                            (32'h3002100c)
`define SOC_SHA512_ACC_CSR_DLEN                                                                     (32'h30021010)
`define SOC_SHA512_ACC_CSR_DATAIN                                                                   (32'h30021014)
`define SOC_SHA512_ACC_CSR_EXECUTE                                                                  (32'h30021018)
`define SOC_SHA512_ACC_CSR_STATUS                                                                   (32'h3002101c)
`define SOC_SHA512_ACC_CSR_DIGEST_0                                                                 (32'h30021020)
`define SOC_SHA512_ACC_CSR_DIGEST_1                                                                 (32'h30021024)
`define SOC_SHA512_ACC_CSR_DIGEST_2                                                                 (32'h30021028)
`define SOC_SHA512_ACC_CSR_DIGEST_3                                                                 (32'h3002102c)
`define SOC_SHA512_ACC_CSR_DIGEST_4                                                                 (32'h30021030)
`define SOC_SHA512_ACC_CSR_DIGEST_5                                                                 (32'h30021034)
`define SOC_SHA512_ACC_CSR_DIGEST_6                                                                 (32'h30021038)
`define SOC_SHA512_ACC_CSR_DIGEST_7                                                                 (32'h3002103c)
`define SOC_SHA512_ACC_CSR_DIGEST_8                                                                 (32'h30021040)
`define SOC_SHA512_ACC_CSR_DIGEST_9                                                                 (32'h30021044)
`define SOC_SHA512_ACC_CSR_DIGEST_10                                                                (32'h30021048)
`define SOC_SHA512_ACC_CSR_DIGEST_11                                                                (32'h3002104c)
`define SOC_SHA512_ACC_CSR_DIGEST_12                                                                (32'h30021050)
`define SOC_SHA512_ACC_CSR_DIGEST_13                                                                (32'h30021054)
`define SOC_SHA512_ACC_CSR_DIGEST_14                                                                (32'h30021058)
`define SOC_SHA512_ACC_CSR_DIGEST_15                                                                (32'h3002105c)
`define SOC_SHA512_ACC_CSR_CONTROL                                                                  (32'h30021060)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_START                                                      (32'h30021800)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                           (32'h30021800)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                            (32'h30021804)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                            (32'h30021808)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                        (32'h3002180c)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                        (32'h30021810)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                      (32'h30021814)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                      (32'h30021818)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                          (32'h3002181c)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                          (32'h30021820)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                        (32'h30021900)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                        (32'h30021904)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                        (32'h30021908)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                        (32'h3002190c)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                (32'h30021980)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                   (32'h30021a00)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                   (32'h30021a04)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                   (32'h30021a08)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                   (32'h30021a0c)
`define SOC_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                           (32'h30021a10)
`define SOC_SOC_IFC_REG_BASE_ADDR                                                                   (32'h30030000)
`define SOC_SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                        (32'h30030000)
`define SOC_SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                    (32'h30030004)
`define SOC_SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                        (32'h30030008)
`define SOC_SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                    (32'h3003000c)
`define SOC_SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                          (32'h30030010)
`define SOC_SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                          (32'h30030014)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                              (32'h30030018)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                              (32'h3003001c)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                              (32'h30030020)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                              (32'h30030024)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                              (32'h30030028)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                              (32'h3003002c)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                              (32'h30030030)
`define SOC_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                              (32'h30030034)
`define SOC_SOC_IFC_REG_CPTRA_BOOT_STATUS                                                           (32'h30030038)
`define SOC_SOC_IFC_REG_CPTRA_FLOW_STATUS                                                           (32'h3003003c)
`define SOC_SOC_IFC_REG_CPTRA_RESET_REASON                                                          (32'h30030040)
`define SOC_SOC_IFC_REG_CPTRA_SECURITY_STATE                                                        (32'h30030044)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_0                                                 (32'h30030048)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_1                                                 (32'h3003004c)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_2                                                 (32'h30030050)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_3                                                 (32'h30030054)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_4                                                 (32'h30030058)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_0                                                  (32'h3003005c)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_1                                                  (32'h30030060)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_2                                                  (32'h30030064)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_3                                                  (32'h30030068)
`define SOC_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_4                                                  (32'h3003006c)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_VALID_AXI_USER                                                   (32'h30030070)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_AXI_USER_LOCK                                                    (32'h30030074)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                           (32'h30030078)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                           (32'h3003007c)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                           (32'h30030080)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                           (32'h30030084)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                           (32'h30030088)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                           (32'h3003008c)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                           (32'h30030090)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                           (32'h30030094)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                           (32'h30030098)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                           (32'h3003009c)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                          (32'h300300a0)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                          (32'h300300a4)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_CTRL                                                             (32'h300300a8)
`define SOC_SOC_IFC_REG_CPTRA_TRNG_STATUS                                                           (32'h300300ac)
`define SOC_SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                          (32'h300300b0)
`define SOC_SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                          (32'h300300b4)
`define SOC_SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                            (32'h300300b8)
`define SOC_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                 (32'h300300bc)
`define SOC_SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                         (32'h300300c0)
`define SOC_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                 (32'h300300c4)
`define SOC_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                 (32'h300300c8)
`define SOC_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                (32'h300300cc)
`define SOC_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                (32'h300300d0)
`define SOC_SOC_IFC_REG_CPTRA_HW_REV_ID                                                             (32'h300300d4)
`define SOC_SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                           (32'h300300d8)
`define SOC_SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                           (32'h300300dc)
`define SOC_SOC_IFC_REG_CPTRA_HW_CONFIG                                                             (32'h300300e0)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER1_EN                                                         (32'h300300e4)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL                                                       (32'h300300e8)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                                           (32'h300300ec)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                                           (32'h300300f0)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER2_EN                                                         (32'h300300f4)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL                                                       (32'h300300f8)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                                           (32'h300300fc)
`define SOC_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                                           (32'h30030100)
`define SOC_SOC_IFC_REG_CPTRA_WDT_STATUS                                                            (32'h30030104)
`define SOC_SOC_IFC_REG_CPTRA_FUSE_VALID_AXI_USER                                                   (32'h30030108)
`define SOC_SOC_IFC_REG_CPTRA_FUSE_AXI_USER_LOCK                                                    (32'h3003010c)
`define SOC_SOC_IFC_REG_CPTRA_WDT_CFG_0                                                             (32'h30030110)
`define SOC_SOC_IFC_REG_CPTRA_WDT_CFG_1                                                             (32'h30030114)
`define SOC_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                                                (32'h30030118)
`define SOC_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                                                (32'h3003011c)
`define SOC_SOC_IFC_REG_CPTRA_RSVD_REG_0                                                            (32'h30030120)
`define SOC_SOC_IFC_REG_CPTRA_RSVD_REG_1                                                            (32'h30030124)
`define SOC_SOC_IFC_REG_CPTRA_HW_CAPABILITIES                                                       (32'h30030128)
`define SOC_SOC_IFC_REG_CPTRA_FW_CAPABILITIES                                                       (32'h3003012c)
`define SOC_SOC_IFC_REG_CPTRA_CAP_LOCK                                                              (32'h30030130)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_0                                                       (32'h30030140)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_1                                                       (32'h30030144)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_2                                                       (32'h30030148)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_3                                                       (32'h3003014c)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_4                                                       (32'h30030150)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_5                                                       (32'h30030154)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_6                                                       (32'h30030158)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_7                                                       (32'h3003015c)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_8                                                       (32'h30030160)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_9                                                       (32'h30030164)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_10                                                      (32'h30030168)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_11                                                      (32'h3003016c)
`define SOC_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_LOCK                                                    (32'h30030170)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_0                                                             (32'h30030200)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_1                                                             (32'h30030204)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_2                                                             (32'h30030208)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_3                                                             (32'h3003020c)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_4                                                             (32'h30030210)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_5                                                             (32'h30030214)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_6                                                             (32'h30030218)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_7                                                             (32'h3003021c)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_8                                                             (32'h30030220)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_9                                                             (32'h30030224)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_10                                                            (32'h30030228)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_11                                                            (32'h3003022c)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_12                                                            (32'h30030230)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_13                                                            (32'h30030234)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_14                                                            (32'h30030238)
`define SOC_SOC_IFC_REG_FUSE_UDS_SEED_15                                                            (32'h3003023c)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                        (32'h30030240)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                        (32'h30030244)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                        (32'h30030248)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                        (32'h3003024c)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                        (32'h30030250)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                        (32'h30030254)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                        (32'h30030258)
`define SOC_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                        (32'h3003025c)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_0                                                       (32'h30030260)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_1                                                       (32'h30030264)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_2                                                       (32'h30030268)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_3                                                       (32'h3003026c)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_4                                                       (32'h30030270)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_5                                                       (32'h30030274)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_6                                                       (32'h30030278)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_7                                                       (32'h3003027c)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_8                                                       (32'h30030280)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_9                                                       (32'h30030284)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_10                                                      (32'h30030288)
`define SOC_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_11                                                      (32'h3003028c)
`define SOC_SOC_IFC_REG_FUSE_ECC_REVOCATION                                                         (32'h30030290)
`define SOC_SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                   (32'h300302b4)
`define SOC_SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                          (32'h300302b8)
`define SOC_SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                          (32'h300302bc)
`define SOC_SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                          (32'h300302c0)
`define SOC_SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                          (32'h300302c4)
`define SOC_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                  (32'h300302c8)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                     (32'h300302cc)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                     (32'h300302d0)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                     (32'h300302d4)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                     (32'h300302d8)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                     (32'h300302dc)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                     (32'h300302e0)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                     (32'h300302e4)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                     (32'h300302e8)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                     (32'h300302ec)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                     (32'h300302f0)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                    (32'h300302f4)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                    (32'h300302f8)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                    (32'h300302fc)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                    (32'h30030300)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                    (32'h30030304)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                    (32'h30030308)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                    (32'h3003030c)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                    (32'h30030310)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                    (32'h30030314)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                    (32'h30030318)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                    (32'h3003031c)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                    (32'h30030320)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                    (32'h30030324)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                    (32'h30030328)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                  (32'h3003032c)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                  (32'h30030330)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                  (32'h30030334)
`define SOC_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                  (32'h30030338)
`define SOC_SOC_IFC_REG_FUSE_LMS_REVOCATION                                                         (32'h30030340)
`define SOC_SOC_IFC_REG_FUSE_MLDSA_REVOCATION                                                       (32'h30030344)
`define SOC_SOC_IFC_REG_FUSE_SOC_STEPPING_ID                                                        (32'h30030348)
`define SOC_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_0                                               (32'h3003034c)
`define SOC_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_1                                               (32'h30030350)
`define SOC_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_2                                               (32'h30030354)
`define SOC_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_3                                               (32'h30030358)
`define SOC_SOC_IFC_REG_FUSE_PQC_KEY_TYPE                                                           (32'h3003035c)
`define SOC_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_0                                                     (32'h30030360)
`define SOC_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_1                                                     (32'h30030364)
`define SOC_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_2                                                     (32'h30030368)
`define SOC_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_3                                                     (32'h3003036c)
`define SOC_SOC_IFC_REG_FUSE_SOC_MANIFEST_MAX_SVN                                                   (32'h30030370)
`define SOC_SOC_IFC_REG_SS_CALIPTRA_BASE_ADDR_L                                                     (32'h30030500)
`define SOC_SOC_IFC_REG_SS_CALIPTRA_BASE_ADDR_H                                                     (32'h30030504)
`define SOC_SOC_IFC_REG_SS_MCI_BASE_ADDR_L                                                          (32'h30030508)
`define SOC_SOC_IFC_REG_SS_MCI_BASE_ADDR_H                                                          (32'h3003050c)
`define SOC_SOC_IFC_REG_SS_RECOVERY_IFC_BASE_ADDR_L                                                 (32'h30030510)
`define SOC_SOC_IFC_REG_SS_RECOVERY_IFC_BASE_ADDR_H                                                 (32'h30030514)
`define SOC_SOC_IFC_REG_SS_OTP_FC_BASE_ADDR_L                                                       (32'h30030518)
`define SOC_SOC_IFC_REG_SS_OTP_FC_BASE_ADDR_H                                                       (32'h3003051c)
`define SOC_SOC_IFC_REG_SS_UDS_SEED_BASE_ADDR_L                                                     (32'h30030520)
`define SOC_SOC_IFC_REG_SS_UDS_SEED_BASE_ADDR_H                                                     (32'h30030524)
`define SOC_SOC_IFC_REG_SS_PROD_DEBUG_UNLOCK_AUTH_PK_HASH_REG_BANK_OFFSET                           (32'h30030528)
`define SOC_SOC_IFC_REG_SS_NUM_OF_PROD_DEBUG_UNLOCK_AUTH_PK_HASHES                                  (32'h3003052c)
`define SOC_SOC_IFC_REG_SS_DEBUG_INTENT                                                             (32'h30030530)
`define SOC_SOC_IFC_REG_SS_CALIPTRA_DMA_AXI_USER                                                    (32'h30030534)
`define SOC_SOC_IFC_REG_SS_STRAP_GENERIC_0                                                          (32'h300305a0)
`define SOC_SOC_IFC_REG_SS_STRAP_GENERIC_1                                                          (32'h300305a4)
`define SOC_SOC_IFC_REG_SS_STRAP_GENERIC_2                                                          (32'h300305a8)
`define SOC_SOC_IFC_REG_SS_STRAP_GENERIC_3                                                          (32'h300305ac)
`define SOC_SOC_IFC_REG_SS_DBG_MANUF_SERVICE_REG_REQ                                                (32'h300305c0)
`define SOC_SOC_IFC_REG_SS_DBG_MANUF_SERVICE_REG_RSP                                                (32'h300305c4)
`define SOC_SOC_IFC_REG_SS_SOC_DBG_UNLOCK_LEVEL_0                                                   (32'h300305c8)
`define SOC_SOC_IFC_REG_SS_SOC_DBG_UNLOCK_LEVEL_1                                                   (32'h300305cc)
`define SOC_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_0                                                   (32'h300305d0)
`define SOC_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_1                                                   (32'h300305d4)
`define SOC_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_2                                                   (32'h300305d8)
`define SOC_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_3                                                   (32'h300305dc)


`endif