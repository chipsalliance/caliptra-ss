// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef MCI_TOP_DEFINES_HEADER
`define MCI_TOP_DEFINES_HEADER


`define MCI_TOP_BASE_ADDR                                                                           (32'h0)
`define MCI_TOP_MCI_REG_BASE_ADDR                                                                   (32'h0)
`define MCI_TOP_MCI_REG_HW_CAPABILITIES                                                             (32'h0)
`define MCI_TOP_MCI_REG_FW_CAPABILITIES                                                             (32'h4)
`define MCI_TOP_MCI_REG_CAP_LOCK                                                                    (32'h8)
`define MCI_TOP_MCI_REG_HW_REV_ID                                                                   (32'hc)
`define MCI_TOP_MCI_REG_FW_REV_ID_0                                                                 (32'h10)
`define MCI_TOP_MCI_REG_FW_REV_ID_1                                                                 (32'h14)
`define MCI_TOP_MCI_REG_HW_CONFIG0                                                                  (32'h18)
`define MCI_TOP_MCI_REG_HW_CONFIG1                                                                  (32'h1c)
`define MCI_TOP_MCI_REG_FW_FLOW_STATUS                                                              (32'h20)
`define MCI_TOP_MCI_REG_HW_FLOW_STATUS                                                              (32'h24)
`define MCI_TOP_MCI_REG_RESET_REASON                                                                (32'h28)
`define MCI_TOP_MCI_REG_RESET_STATUS                                                                (32'h2c)
`define MCI_TOP_MCI_REG_SECURITY_STATE                                                              (32'h30)
`define MCI_TOP_MCI_REG_HW_ERROR_FATAL                                                              (32'h40)
`define MCI_TOP_MCI_REG_AGG_ERROR_FATAL                                                             (32'h44)
`define MCI_TOP_MCI_REG_HW_ERROR_NON_FATAL                                                          (32'h48)
`define MCI_TOP_MCI_REG_AGG_ERROR_NON_FATAL                                                         (32'h4c)
`define MCI_TOP_MCI_REG_FW_ERROR_FATAL                                                              (32'h50)
`define MCI_TOP_MCI_REG_FW_ERROR_NON_FATAL                                                          (32'h54)
`define MCI_TOP_MCI_REG_HW_ERROR_ENC                                                                (32'h58)
`define MCI_TOP_MCI_REG_FW_ERROR_ENC                                                                (32'h5c)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_0                                                    (32'h60)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_1                                                    (32'h64)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_2                                                    (32'h68)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_3                                                    (32'h6c)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_4                                                    (32'h70)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_5                                                    (32'h74)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_6                                                    (32'h78)
`define MCI_TOP_MCI_REG_FW_EXTENDED_ERROR_INFO_7                                                    (32'h7c)
`define MCI_TOP_MCI_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                (32'h80)
`define MCI_TOP_MCI_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                            (32'h84)
`define MCI_TOP_MCI_REG_INTERNAL_AGG_ERROR_FATAL_MASK                                               (32'h88)
`define MCI_TOP_MCI_REG_INTERNAL_AGG_ERROR_NON_FATAL_MASK                                           (32'h8c)
`define MCI_TOP_MCI_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                (32'h90)
`define MCI_TOP_MCI_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                            (32'h94)
`define MCI_TOP_MCI_REG_WDT_TIMER1_EN                                                               (32'ha0)
`define MCI_TOP_MCI_REG_WDT_TIMER1_CTRL                                                             (32'ha4)
`define MCI_TOP_MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_0                                                 (32'ha8)
`define MCI_TOP_MCI_REG_WDT_TIMER1_TIMEOUT_PERIOD_1                                                 (32'hac)
`define MCI_TOP_MCI_REG_WDT_TIMER2_EN                                                               (32'hb0)
`define MCI_TOP_MCI_REG_WDT_TIMER2_CTRL                                                             (32'hb4)
`define MCI_TOP_MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_0                                                 (32'hb8)
`define MCI_TOP_MCI_REG_WDT_TIMER2_TIMEOUT_PERIOD_1                                                 (32'hbc)
`define MCI_TOP_MCI_REG_WDT_STATUS                                                                  (32'hc0)
`define MCI_TOP_MCI_REG_WDT_CFG_0                                                                   (32'hd0)
`define MCI_TOP_MCI_REG_WDT_CFG_1                                                                   (32'hd4)
`define MCI_TOP_MCI_REG_MCU_TIMER_CONFIG                                                            (32'he0)
`define MCI_TOP_MCI_REG_MCU_RV_MTIME_L                                                              (32'he4)
`define MCI_TOP_MCI_REG_MCU_RV_MTIME_H                                                              (32'he8)
`define MCI_TOP_MCI_REG_MCU_RV_MTIMECMP_L                                                           (32'hec)
`define MCI_TOP_MCI_REG_MCU_RV_MTIMECMP_H                                                           (32'hf0)
`define MCI_TOP_MCI_REG_RESET_REQUEST                                                               (32'h100)
`define MCI_TOP_MCI_REG_MCI_BOOTFSM_GO                                                              (32'h104)
`define MCI_TOP_MCI_REG_CPTRA_BOOT_GO                                                               (32'h108)
`define MCI_TOP_MCI_REG_FW_SRAM_EXEC_REGION_SIZE                                                    (32'h10c)
`define MCI_TOP_MCI_REG_MCU_NMI_VECTOR                                                              (32'h110)
`define MCI_TOP_MCI_REG_MCU_RESET_VECTOR                                                            (32'h114)
`define MCI_TOP_MCI_REG_MBOX0_VALID_AXI_USER_0                                                      (32'h180)
`define MCI_TOP_MCI_REG_MBOX0_VALID_AXI_USER_1                                                      (32'h184)
`define MCI_TOP_MCI_REG_MBOX0_VALID_AXI_USER_2                                                      (32'h188)
`define MCI_TOP_MCI_REG_MBOX0_VALID_AXI_USER_3                                                      (32'h18c)
`define MCI_TOP_MCI_REG_MBOX0_VALID_AXI_USER_4                                                      (32'h190)
`define MCI_TOP_MCI_REG_MBOX0_AXI_USER_LOCK_0                                                       (32'h1a0)
`define MCI_TOP_MCI_REG_MBOX0_AXI_USER_LOCK_1                                                       (32'h1a4)
`define MCI_TOP_MCI_REG_MBOX0_AXI_USER_LOCK_2                                                       (32'h1a8)
`define MCI_TOP_MCI_REG_MBOX0_AXI_USER_LOCK_3                                                       (32'h1ac)
`define MCI_TOP_MCI_REG_MBOX0_AXI_USER_LOCK_4                                                       (32'h1b0)
`define MCI_TOP_MCI_REG_MBOX1_VALID_AXI_USER_0                                                      (32'h1c0)
`define MCI_TOP_MCI_REG_MBOX1_VALID_AXI_USER_1                                                      (32'h1c4)
`define MCI_TOP_MCI_REG_MBOX1_VALID_AXI_USER_2                                                      (32'h1c8)
`define MCI_TOP_MCI_REG_MBOX1_VALID_AXI_USER_3                                                      (32'h1cc)
`define MCI_TOP_MCI_REG_MBOX1_VALID_AXI_USER_4                                                      (32'h1d0)
`define MCI_TOP_MCI_REG_MBOX1_AXI_USER_LOCK_0                                                       (32'h1e0)
`define MCI_TOP_MCI_REG_MBOX1_AXI_USER_LOCK_1                                                       (32'h1e4)
`define MCI_TOP_MCI_REG_MBOX1_AXI_USER_LOCK_2                                                       (32'h1e8)
`define MCI_TOP_MCI_REG_MBOX1_AXI_USER_LOCK_3                                                       (32'h1ec)
`define MCI_TOP_MCI_REG_MBOX1_AXI_USER_LOCK_4                                                       (32'h1f0)
`define MCI_TOP_MCI_REG_SOC_DFT_EN_0                                                                (32'h300)
`define MCI_TOP_MCI_REG_SOC_DFT_EN_1                                                                (32'h304)
`define MCI_TOP_MCI_REG_SOC_HW_DEBUG_EN_0                                                           (32'h308)
`define MCI_TOP_MCI_REG_SOC_HW_DEBUG_EN_1                                                           (32'h30c)
`define MCI_TOP_MCI_REG_SOC_PROD_DEBUG_STATE_0                                                      (32'h310)
`define MCI_TOP_MCI_REG_SOC_PROD_DEBUG_STATE_1                                                      (32'h314)
`define MCI_TOP_MCI_REG_FC_FIPS_ZEROZATION                                                          (32'h318)
`define MCI_TOP_MCI_REG_GENERIC_INPUT_WIRES_0                                                       (32'h400)
`define MCI_TOP_MCI_REG_GENERIC_INPUT_WIRES_1                                                       (32'h404)
`define MCI_TOP_MCI_REG_GENERIC_OUTPUT_WIRES_0                                                      (32'h408)
`define MCI_TOP_MCI_REG_GENERIC_OUTPUT_WIRES_1                                                      (32'h40c)
`define MCI_TOP_MCI_REG_DEBUG_IN                                                                    (32'h410)
`define MCI_TOP_MCI_REG_DEBUG_OUT                                                                   (32'h414)
`define MCI_TOP_MCI_REG_SS_DEBUG_INTENT                                                             (32'h418)
`define MCI_TOP_MCI_REG_SS_CONFIG_DONE_STICKY                                                       (32'h440)
`define MCI_TOP_MCI_REG_SS_CONFIG_DONE                                                              (32'h444)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_0                                           (32'h480)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_1                                           (32'h484)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_2                                           (32'h488)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_3                                           (32'h48c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_4                                           (32'h490)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_5                                           (32'h494)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_6                                           (32'h498)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_7                                           (32'h49c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_8                                           (32'h4a0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_9                                           (32'h4a4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_10                                          (32'h4a8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_0_11                                          (32'h4ac)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_0                                           (32'h4b0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_1                                           (32'h4b4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_2                                           (32'h4b8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_3                                           (32'h4bc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_4                                           (32'h4c0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_5                                           (32'h4c4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_6                                           (32'h4c8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_7                                           (32'h4cc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_8                                           (32'h4d0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_9                                           (32'h4d4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_10                                          (32'h4d8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_1_11                                          (32'h4dc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_0                                           (32'h4e0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_1                                           (32'h4e4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_2                                           (32'h4e8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_3                                           (32'h4ec)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_4                                           (32'h4f0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_5                                           (32'h4f4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_6                                           (32'h4f8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_7                                           (32'h4fc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_8                                           (32'h500)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_9                                           (32'h504)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_10                                          (32'h508)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_2_11                                          (32'h50c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_0                                           (32'h510)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_1                                           (32'h514)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_2                                           (32'h518)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_3                                           (32'h51c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_4                                           (32'h520)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_5                                           (32'h524)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_6                                           (32'h528)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_7                                           (32'h52c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_8                                           (32'h530)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_9                                           (32'h534)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_10                                          (32'h538)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_3_11                                          (32'h53c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_0                                           (32'h540)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_1                                           (32'h544)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_2                                           (32'h548)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_3                                           (32'h54c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_4                                           (32'h550)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_5                                           (32'h554)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_6                                           (32'h558)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_7                                           (32'h55c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_8                                           (32'h560)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_9                                           (32'h564)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_10                                          (32'h568)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_4_11                                          (32'h56c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_0                                           (32'h570)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_1                                           (32'h574)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_2                                           (32'h578)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_3                                           (32'h57c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_4                                           (32'h580)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_5                                           (32'h584)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_6                                           (32'h588)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_7                                           (32'h58c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_8                                           (32'h590)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_9                                           (32'h594)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_10                                          (32'h598)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_5_11                                          (32'h59c)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_0                                           (32'h5a0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_1                                           (32'h5a4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_2                                           (32'h5a8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_3                                           (32'h5ac)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_4                                           (32'h5b0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_5                                           (32'h5b4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_6                                           (32'h5b8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_7                                           (32'h5bc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_8                                           (32'h5c0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_9                                           (32'h5c4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_10                                          (32'h5c8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_6_11                                          (32'h5cc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_0                                           (32'h5d0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_1                                           (32'h5d4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_2                                           (32'h5d8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_3                                           (32'h5dc)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_4                                           (32'h5e0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_5                                           (32'h5e4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_6                                           (32'h5e8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_7                                           (32'h5ec)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_8                                           (32'h5f0)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_9                                           (32'h5f4)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_10                                          (32'h5f8)
`define MCI_TOP_MCI_REG_PROD_DEBUG_UNLOCK_PK_HASH_REG_7_11                                          (32'h5fc)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_START                                                         (32'h1000)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h1000)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_EN_R                                              (32'h1004)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_EN_R                                              (32'h1008)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_EN_R                                              (32'h100c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_EN_R                                              (32'h1010)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h1014)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h1018)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR0_INTERNAL_INTR_R                                        (32'h101c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR1_INTERNAL_INTR_R                                        (32'h1020)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTERNAL_INTR_R                                        (32'h1024)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTERNAL_INTR_R                                        (32'h1028)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR0_INTR_TRIG_R                                            (32'h102c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR1_INTR_TRIG_R                                            (32'h1030)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF0_INTR_TRIG_R                                            (32'h1034)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF1_INTR_TRIG_R                                            (32'h1038)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                   (32'h1100)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_INV_DEV_INTR_COUNT_R                              (32'h1104)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_INV_DEV_INTR_COUNT_R                              (32'h1108)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_CMD_FAIL_INTR_COUNT_R                             (32'h110c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_CMD_FAIL_INTR_COUNT_R                             (32'h1110)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_ECC_UNC_INTR_COUNT_R                              (32'h1114)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_ECC_UNC_INTR_COUNT_R                              (32'h1118)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MCU_SRAM_DMI_AXI_COLLISION_INTR_COUNT_R                 (32'h111c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                         (32'h1120)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                         (32'h1124)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_R                           (32'h1128)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_R                           (32'h112c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_R                           (32'h1130)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_R                           (32'h1134)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_R                           (32'h1138)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_R                           (32'h113c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_R                           (32'h1140)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_R                           (32'h1144)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_R                           (32'h1148)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_R                           (32'h114c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_R                          (32'h1150)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_R                          (32'h1154)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_R                          (32'h1158)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_R                          (32'h115c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_R                          (32'h1160)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_R                          (32'h1164)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_R                          (32'h1168)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_R                          (32'h116c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_R                          (32'h1170)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_R                          (32'h1174)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_R                          (32'h1178)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_R                          (32'h117c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_R                          (32'h1180)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_R                          (32'h1184)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_R                          (32'h1188)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_R                          (32'h118c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_R                          (32'h1190)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_R                          (32'h1194)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_R                          (32'h1198)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_R                          (32'h119c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_R                          (32'h11a0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_R                          (32'h11a4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_R                           (32'h1200)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MCU_RESET_REQ_INTR_COUNT_R                        (32'h1204)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_R                              (32'h1208)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_R                       (32'h120c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_R                       (32'h1210)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_R                       (32'h1214)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_R                       (32'h1218)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_R                       (32'h121c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_R                       (32'h1220)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_R                       (32'h1224)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_R                       (32'h1228)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_R                       (32'h122c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_R                       (32'h1230)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_R                      (32'h1234)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_R                      (32'h1238)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_R                      (32'h123c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_R                      (32'h1240)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_R                      (32'h1244)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_R                      (32'h1248)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_R                      (32'h124c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_R                      (32'h1250)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_R                      (32'h1254)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_R                      (32'h1258)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_R                      (32'h125c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_R                      (32'h1260)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_R                      (32'h1264)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_R                      (32'h1268)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_R                      (32'h126c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_R                      (32'h1270)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_R                      (32'h1274)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_R                      (32'h1278)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_R                      (32'h127c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_R                      (32'h1280)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_R                      (32'h1284)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_R                      (32'h1288)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_CMD_AVAIL_INTR_COUNT_R                            (32'h128c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_CMD_AVAIL_INTR_COUNT_R                            (32'h1290)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MBOX_CMD_AVAIL_INTR_COUNT_R                       (32'h1294)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_ECC_COR_INTR_COUNT_R                              (32'h1298)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_ECC_COR_INTR_COUNT_R                              (32'h129c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                               (32'h12a0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_R                                  (32'h12a4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_SOC_REQ_LOCK_INTR_COUNT_R                         (32'h12a8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_SOC_REQ_LOCK_INTR_COUNT_R                         (32'h12ac)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                              (32'h1300)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_INV_DEV_INTR_COUNT_INCR_R                         (32'h1304)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_INV_DEV_INTR_COUNT_INCR_R                         (32'h1308)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_CMD_FAIL_INTR_COUNT_INCR_R                        (32'h130c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_CMD_FAIL_INTR_COUNT_INCR_R                        (32'h1310)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX0_ECC_UNC_INTR_COUNT_INCR_R                         (32'h1314)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MBOX1_ECC_UNC_INTR_COUNT_INCR_R                         (32'h1318)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                    (32'h131c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                    (32'h1320)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_MCU_SRAM_DMI_AXI_COLLISION_INTR_COUNT_INCR_R            (32'h1324)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL0_INTR_COUNT_INCR_R                      (32'h1328)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL1_INTR_COUNT_INCR_R                      (32'h132c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL2_INTR_COUNT_INCR_R                      (32'h1330)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL3_INTR_COUNT_INCR_R                      (32'h1334)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL4_INTR_COUNT_INCR_R                      (32'h1338)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL5_INTR_COUNT_INCR_R                      (32'h133c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL6_INTR_COUNT_INCR_R                      (32'h1340)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL7_INTR_COUNT_INCR_R                      (32'h1344)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL8_INTR_COUNT_INCR_R                      (32'h1348)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL9_INTR_COUNT_INCR_R                      (32'h134c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL10_INTR_COUNT_INCR_R                     (32'h1350)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL11_INTR_COUNT_INCR_R                     (32'h1354)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL12_INTR_COUNT_INCR_R                     (32'h1358)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL13_INTR_COUNT_INCR_R                     (32'h135c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL14_INTR_COUNT_INCR_R                     (32'h1360)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL15_INTR_COUNT_INCR_R                     (32'h1364)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL16_INTR_COUNT_INCR_R                     (32'h1368)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL17_INTR_COUNT_INCR_R                     (32'h136c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL18_INTR_COUNT_INCR_R                     (32'h1370)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL19_INTR_COUNT_INCR_R                     (32'h1374)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL20_INTR_COUNT_INCR_R                     (32'h1378)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL21_INTR_COUNT_INCR_R                     (32'h137c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL22_INTR_COUNT_INCR_R                     (32'h1380)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL23_INTR_COUNT_INCR_R                     (32'h1384)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL24_INTR_COUNT_INCR_R                     (32'h1388)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL25_INTR_COUNT_INCR_R                     (32'h138c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL26_INTR_COUNT_INCR_R                     (32'h1390)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL27_INTR_COUNT_INCR_R                     (32'h1394)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL28_INTR_COUNT_INCR_R                     (32'h1398)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL29_INTR_COUNT_INCR_R                     (32'h139c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL30_INTR_COUNT_INCR_R                     (32'h13a0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_ERROR_AGG_ERROR_FATAL31_INTR_COUNT_INCR_R                     (32'h13a4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MCU_SRAM_ECC_COR_INTR_COUNT_INCR_R                      (32'h13a8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MCU_RESET_REQ_INTR_COUNT_INCR_R                   (32'h13ac)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R                         (32'h13b0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL0_INTR_COUNT_INCR_R                  (32'h13b4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL1_INTR_COUNT_INCR_R                  (32'h13b8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL2_INTR_COUNT_INCR_R                  (32'h13bc)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL3_INTR_COUNT_INCR_R                  (32'h13c0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL4_INTR_COUNT_INCR_R                  (32'h13c4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL5_INTR_COUNT_INCR_R                  (32'h13c8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL6_INTR_COUNT_INCR_R                  (32'h13cc)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL7_INTR_COUNT_INCR_R                  (32'h13d0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL8_INTR_COUNT_INCR_R                  (32'h13d4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL9_INTR_COUNT_INCR_R                  (32'h13d8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL10_INTR_COUNT_INCR_R                 (32'h13dc)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL11_INTR_COUNT_INCR_R                 (32'h13e0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL12_INTR_COUNT_INCR_R                 (32'h13e4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL13_INTR_COUNT_INCR_R                 (32'h13e8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL14_INTR_COUNT_INCR_R                 (32'h13ec)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL15_INTR_COUNT_INCR_R                 (32'h13f0)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL16_INTR_COUNT_INCR_R                 (32'h13f4)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL17_INTR_COUNT_INCR_R                 (32'h13f8)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL18_INTR_COUNT_INCR_R                 (32'h13fc)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL19_INTR_COUNT_INCR_R                 (32'h1400)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL20_INTR_COUNT_INCR_R                 (32'h1404)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL21_INTR_COUNT_INCR_R                 (32'h1408)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL22_INTR_COUNT_INCR_R                 (32'h140c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL23_INTR_COUNT_INCR_R                 (32'h1410)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL24_INTR_COUNT_INCR_R                 (32'h1414)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL25_INTR_COUNT_INCR_R                 (32'h1418)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL26_INTR_COUNT_INCR_R                 (32'h141c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL27_INTR_COUNT_INCR_R                 (32'h1420)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL28_INTR_COUNT_INCR_R                 (32'h1424)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL29_INTR_COUNT_INCR_R                 (32'h1428)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL30_INTR_COUNT_INCR_R                 (32'h142c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_AGG_ERROR_NON_FATAL31_INTR_COUNT_INCR_R                 (32'h1430)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_CMD_AVAIL_INTR_COUNT_INCR_R                       (32'h1434)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_CMD_AVAIL_INTR_COUNT_INCR_R                       (32'h1438)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_CPTRA_MBOX_CMD_AVAIL_INTR_COUNT_INCR_R                  (32'h143c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_ECC_COR_INTR_COUNT_INCR_R                         (32'h1440)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_ECC_COR_INTR_COUNT_INCR_R                         (32'h1444)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                          (32'h1448)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R                             (32'h144c)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX0_SOC_REQ_LOCK_INTR_COUNT_INCR_R                    (32'h1450)
`define MCI_TOP_MCI_REG_INTR_BLOCK_RF_NOTIF_MBOX1_SOC_REQ_LOCK_INTR_COUNT_INCR_R                    (32'h1454)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_BASE_ADDR                                                      (32'h10000)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_STATUS                                                         (32'h10000)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_CONFIG                                                         (32'h10004)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_DATA                                                           (32'h10008)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_WRITE_PTR                                                      (32'h1000c)
`define MCI_TOP_MCU_TRACE_BUFFER_CSR_READ_PTR                                                       (32'h10010)
`define MCI_TOP_MBOX0_CSR_BASE_ADDR                                                                 (32'h80000)
`define MCI_TOP_MBOX0_CSR_MBOX_LOCK                                                                 (32'h80000)
`define MCI_TOP_MBOX0_CSR_MBOX_USER                                                                 (32'h80004)
`define MCI_TOP_MBOX0_CSR_MBOX_CMD                                                                  (32'h80008)
`define MCI_TOP_MBOX0_CSR_MBOX_DLEN                                                                 (32'h8000c)
`define MCI_TOP_MBOX0_CSR_MBOX_DATAIN                                                               (32'h80010)
`define MCI_TOP_MBOX0_CSR_MBOX_DATAOUT                                                              (32'h80014)
`define MCI_TOP_MBOX0_CSR_MBOX_EXECUTE                                                              (32'h80018)
`define MCI_TOP_MBOX0_CSR_MBOX_STATUS                                                               (32'h8001c)
`define MCI_TOP_MBOX0_CSR_MBOX_UNLOCK                                                               (32'h80020)
`define MCI_TOP_MBOX0_CSR_TAP_MODE                                                                  (32'h80024)
`define MCI_TOP_MBOX1_CSR_BASE_ADDR                                                                 (32'h90000)
`define MCI_TOP_MBOX1_CSR_MBOX_LOCK                                                                 (32'h90000)
`define MCI_TOP_MBOX1_CSR_MBOX_USER                                                                 (32'h90004)
`define MCI_TOP_MBOX1_CSR_MBOX_CMD                                                                  (32'h90008)
`define MCI_TOP_MBOX1_CSR_MBOX_DLEN                                                                 (32'h9000c)
`define MCI_TOP_MBOX1_CSR_MBOX_DATAIN                                                               (32'h90010)
`define MCI_TOP_MBOX1_CSR_MBOX_DATAOUT                                                              (32'h90014)
`define MCI_TOP_MBOX1_CSR_MBOX_EXECUTE                                                              (32'h90018)
`define MCI_TOP_MBOX1_CSR_MBOX_STATUS                                                               (32'h9001c)
`define MCI_TOP_MBOX1_CSR_MBOX_UNLOCK                                                               (32'h90020)
`define MCI_TOP_MBOX1_CSR_TAP_MODE                                                                  (32'h90024)
`define MCI_TOP_MCU_SRAM_BASE_ADDR                                                                  (32'h200000)
`define MCI_TOP_MCU_SRAM_END_ADDR                                                                   (32'h3fffff)


`endif