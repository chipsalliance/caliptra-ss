
`ifndef CPTRA_SS_INCLUDES_SVH
`define CPTRA_SS_INCLUDES_SVH


parameter CPTRA_SS_MCU_USER_WIDTH               = 32;
parameter CPTRA_SS_STRAP_CLPTRA_CORE_AXI_USER   = 32'hFFFF_FFFF;
parameter CPTRA_SS_STRAP_MCU_LSU_AXI_USER       = 32'h1;

`endif // CPTRA_SS_INCLUDES_SVH