// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//



`include "caliptra_prim_assert.sv"

module otp_ctrl_prim_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output otp_ctrl_reg_pkg::otp_ctrl_prim_reg2hw_t reg2hw, // Write
  input  otp_ctrl_reg_pkg::otp_ctrl_prim_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o
);

  import otp_ctrl_reg_pkg::* ;

  localparam int AW = 5;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [7:0] reg_we_check;
  caliptra_prim_reg_we_check #(
    .OneHotWidth(8)
  ) u_caliptra_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(caliptra_prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = addrmiss | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic csr0_we;
  logic csr0_field0_qs;
  logic csr0_field0_wd;
  logic csr0_field1_qs;
  logic csr0_field1_wd;
  logic csr0_field2_qs;
  logic csr0_field2_wd;
  logic [9:0] csr0_field3_qs;
  logic [9:0] csr0_field3_wd;
  logic [10:0] csr0_field4_qs;
  logic [10:0] csr0_field4_wd;
  logic csr1_we;
  logic [6:0] csr1_field0_qs;
  logic [6:0] csr1_field0_wd;
  logic csr1_field1_qs;
  logic csr1_field1_wd;
  logic [6:0] csr1_field2_qs;
  logic [6:0] csr1_field2_wd;
  logic csr1_field3_qs;
  logic csr1_field3_wd;
  logic [15:0] csr1_field4_qs;
  logic [15:0] csr1_field4_wd;
  logic csr2_we;
  logic csr2_qs;
  logic csr2_wd;
  logic csr3_we;
  logic [2:0] csr3_field0_qs;
  logic [2:0] csr3_field0_wd;
  logic [9:0] csr3_field1_qs;
  logic [9:0] csr3_field1_wd;
  logic csr3_field2_qs;
  logic csr3_field2_wd;
  logic csr3_field3_qs;
  logic csr3_field4_qs;
  logic csr3_field5_qs;
  logic csr3_field6_qs;
  logic csr3_field7_qs;
  logic csr3_field8_qs;
  logic csr4_we;
  logic [9:0] csr4_field0_qs;
  logic [9:0] csr4_field0_wd;
  logic csr4_field1_qs;
  logic csr4_field1_wd;
  logic csr4_field2_qs;
  logic csr4_field2_wd;
  logic csr4_field3_qs;
  logic csr4_field3_wd;
  logic csr5_we;
  logic [5:0] csr5_field0_qs;
  logic [5:0] csr5_field0_wd;
  logic [1:0] csr5_field1_qs;
  logic [1:0] csr5_field1_wd;
  logic csr5_field2_qs;
  logic [2:0] csr5_field3_qs;
  logic csr5_field4_qs;
  logic csr5_field5_qs;
  logic [15:0] csr5_field6_qs;
  logic [15:0] csr5_field6_wd;
  logic csr6_we;
  logic [9:0] csr6_field0_qs;
  logic [9:0] csr6_field0_wd;
  logic csr6_field1_qs;
  logic csr6_field1_wd;
  logic csr6_field2_qs;
  logic csr6_field2_wd;
  logic [15:0] csr6_field3_qs;
  logic [15:0] csr6_field3_wd;
  logic [5:0] csr7_field0_qs;
  logic [2:0] csr7_field1_qs;
  logic csr7_field2_qs;
  logic csr7_field3_qs;

  // Register instances
  // R[csr0]: V(False)
  //   F[field0]: 0:0
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr0_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr0_we),
    .wd     (csr0_field0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr0.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr0_field0_qs)
  );

  //   F[field1]: 1:1
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr0_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr0_we),
    .wd     (csr0_field1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr0.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr0_field1_qs)
  );

  //   F[field2]: 2:2
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr0_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr0_we),
    .wd     (csr0_field2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr0.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr0_field2_qs)
  );

  //   F[field3]: 13:4
  caliptra_prim_subreg #(
    .DW      (10),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (10'h0),
    .Mubi    (1'b0)
  ) u_csr0_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr0_we),
    .wd     (csr0_field3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr0.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr0_field3_qs)
  );

  //   F[field4]: 26:16
  caliptra_prim_subreg #(
    .DW      (11),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (11'h0),
    .Mubi    (1'b0)
  ) u_csr0_field4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr0_we),
    .wd     (csr0_field4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr0.field4.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr0_field4_qs)
  );


  // R[csr1]: V(False)
  //   F[field0]: 6:0
  caliptra_prim_subreg #(
    .DW      (7),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (7'h0),
    .Mubi    (1'b0)
  ) u_csr1_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr1_we),
    .wd     (csr1_field0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr1.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr1_field0_qs)
  );

  //   F[field1]: 7:7
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr1_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr1_we),
    .wd     (csr1_field1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr1.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr1_field1_qs)
  );

  //   F[field2]: 14:8
  caliptra_prim_subreg #(
    .DW      (7),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (7'h0),
    .Mubi    (1'b0)
  ) u_csr1_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr1_we),
    .wd     (csr1_field2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr1.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr1_field2_qs)
  );

  //   F[field3]: 15:15
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr1_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr1_we),
    .wd     (csr1_field3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr1.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr1_field3_qs)
  );

  //   F[field4]: 31:16
  caliptra_prim_subreg #(
    .DW      (16),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h0),
    .Mubi    (1'b0)
  ) u_csr1_field4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr1_we),
    .wd     (csr1_field4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr1.field4.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr1_field4_qs)
  );


  // R[csr2]: V(False)
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr2_we),
    .wd     (csr2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr2_qs)
  );


  // R[csr3]: V(False)
  //   F[field0]: 2:0
  caliptra_prim_subreg #(
    .DW      (3),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (3'h0),
    .Mubi    (1'b0)
  ) u_csr3_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr3_we),
    .wd     (csr3_field0_wd),

    // from internal hardware
    .de     (hw2reg.csr3.field0.de),
    .d      (hw2reg.csr3.field0.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field0_qs)
  );

  //   F[field1]: 13:4
  caliptra_prim_subreg #(
    .DW      (10),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (10'h0),
    .Mubi    (1'b0)
  ) u_csr3_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr3_we),
    .wd     (csr3_field1_wd),

    // from internal hardware
    .de     (hw2reg.csr3.field1.de),
    .d      (hw2reg.csr3.field1.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field1_qs)
  );

  //   F[field2]: 16:16
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr3_we),
    .wd     (csr3_field2_wd),

    // from internal hardware
    .de     (hw2reg.csr3.field2.de),
    .d      (hw2reg.csr3.field2.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field2_qs)
  );

  //   F[field3]: 17:17
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field3.de),
    .d      (hw2reg.csr3.field3.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field3_qs)
  );

  //   F[field4]: 18:18
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field4.de),
    .d      (hw2reg.csr3.field4.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field4.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field4_qs)
  );

  //   F[field5]: 19:19
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field5.de),
    .d      (hw2reg.csr3.field5.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field5.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field5_qs)
  );

  //   F[field6]: 20:20
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field6.de),
    .d      (hw2reg.csr3.field6.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field6.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field6_qs)
  );

  //   F[field7]: 21:21
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field7.de),
    .d      (hw2reg.csr3.field7.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field7.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field7_qs)
  );

  //   F[field8]: 22:22
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr3_field8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr3.field8.de),
    .d      (hw2reg.csr3.field8.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr3.field8.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr3_field8_qs)
  );


  // R[csr4]: V(False)
  //   F[field0]: 9:0
  caliptra_prim_subreg #(
    .DW      (10),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (10'h0),
    .Mubi    (1'b0)
  ) u_csr4_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr4_we),
    .wd     (csr4_field0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr4.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr4_field0_qs)
  );

  //   F[field1]: 12:12
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr4_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr4_we),
    .wd     (csr4_field1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr4.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr4_field1_qs)
  );

  //   F[field2]: 13:13
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr4_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr4_we),
    .wd     (csr4_field2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr4.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr4_field2_qs)
  );

  //   F[field3]: 14:14
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr4_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr4_we),
    .wd     (csr4_field3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr4.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr4_field3_qs)
  );


  // R[csr5]: V(False)
  //   F[field0]: 5:0
  caliptra_prim_subreg #(
    .DW      (6),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (6'h0),
    .Mubi    (1'b0)
  ) u_csr5_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr5_we),
    .wd     (csr5_field0_wd),

    // from internal hardware
    .de     (hw2reg.csr5.field0.de),
    .d      (hw2reg.csr5.field0.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field0_qs)
  );

  //   F[field1]: 7:6
  caliptra_prim_subreg #(
    .DW      (2),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (2'h0),
    .Mubi    (1'b0)
  ) u_csr5_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr5_we),
    .wd     (csr5_field1_wd),

    // from internal hardware
    .de     (hw2reg.csr5.field1.de),
    .d      (hw2reg.csr5.field1.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field1_qs)
  );

  //   F[field2]: 8:8
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr5_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr5.field2.de),
    .d      (hw2reg.csr5.field2.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field2_qs)
  );

  //   F[field3]: 11:9
  caliptra_prim_subreg #(
    .DW      (3),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (3'h0),
    .Mubi    (1'b0)
  ) u_csr5_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr5.field3.de),
    .d      (hw2reg.csr5.field3.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field3_qs)
  );

  //   F[field4]: 12:12
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr5_field4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr5.field4.de),
    .d      (hw2reg.csr5.field4.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field4.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field4_qs)
  );

  //   F[field5]: 13:13
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr5_field5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr5.field5.de),
    .d      (hw2reg.csr5.field5.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field5.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field5_qs)
  );

  //   F[field6]: 31:16
  caliptra_prim_subreg #(
    .DW      (16),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h0),
    .Mubi    (1'b0)
  ) u_csr5_field6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr5_we),
    .wd     (csr5_field6_wd),

    // from internal hardware
    .de     (hw2reg.csr5.field6.de),
    .d      (hw2reg.csr5.field6.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr5.field6.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr5_field6_qs)
  );


  // R[csr6]: V(False)
  //   F[field0]: 9:0
  caliptra_prim_subreg #(
    .DW      (10),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (10'h0),
    .Mubi    (1'b0)
  ) u_csr6_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr6_we),
    .wd     (csr6_field0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr6.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr6_field0_qs)
  );

  //   F[field1]: 11:11
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr6_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr6_we),
    .wd     (csr6_field1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr6.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr6_field1_qs)
  );

  //   F[field2]: 12:12
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr6_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr6_we),
    .wd     (csr6_field2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr6.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr6_field2_qs)
  );

  //   F[field3]: 31:16
  caliptra_prim_subreg #(
    .DW      (16),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h0),
    .Mubi    (1'b0)
  ) u_csr6_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (csr6_we),
    .wd     (csr6_field3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr6.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr6_field3_qs)
  );


  // R[csr7]: V(False)
  //   F[field0]: 5:0
  caliptra_prim_subreg #(
    .DW      (6),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (6'h0),
    .Mubi    (1'b0)
  ) u_csr7_field0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr7.field0.de),
    .d      (hw2reg.csr7.field0.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr7.field0.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr7_field0_qs)
  );

  //   F[field1]: 10:8
  caliptra_prim_subreg #(
    .DW      (3),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (3'h0),
    .Mubi    (1'b0)
  ) u_csr7_field1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr7.field1.de),
    .d      (hw2reg.csr7.field1.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr7.field1.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr7_field1_qs)
  );

  //   F[field2]: 14:14
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr7_field2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr7.field2.de),
    .d      (hw2reg.csr7.field2.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr7.field2.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr7_field2_qs)
  );

  //   F[field3]: 15:15
  caliptra_prim_subreg #(
    .DW      (1),
    .SwAccess(caliptra_prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0),
    .Mubi    (1'b0)
  ) u_csr7_field3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.csr7.field3.de),
    .d      (hw2reg.csr7.field3.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.csr7.field3.q),
    .ds     (),

    // to register interface (read)
    .qs     (csr7_field3_qs)
  );



  logic [7:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[0] = (reg_addr == OTP_CTRL_CSR0_OFFSET);
    addr_hit[1] = (reg_addr == OTP_CTRL_CSR1_OFFSET);
    addr_hit[2] = (reg_addr == OTP_CTRL_CSR2_OFFSET);
    addr_hit[3] = (reg_addr == OTP_CTRL_CSR3_OFFSET);
    addr_hit[4] = (reg_addr == OTP_CTRL_CSR4_OFFSET);
    addr_hit[5] = (reg_addr == OTP_CTRL_CSR5_OFFSET);
    addr_hit[6] = (reg_addr == OTP_CTRL_CSR6_OFFSET);
    addr_hit[7] = (reg_addr == OTP_CTRL_CSR7_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[0] & (|(OTP_CTRL_PRIM_PERMIT[0] & ~reg_be))) |
               (addr_hit[1] & (|(OTP_CTRL_PRIM_PERMIT[1] & ~reg_be))) |
               (addr_hit[2] & (|(OTP_CTRL_PRIM_PERMIT[2] & ~reg_be))) |
               (addr_hit[3] & (|(OTP_CTRL_PRIM_PERMIT[3] & ~reg_be))) |
               (addr_hit[4] & (|(OTP_CTRL_PRIM_PERMIT[4] & ~reg_be))) |
               (addr_hit[5] & (|(OTP_CTRL_PRIM_PERMIT[5] & ~reg_be))) |
               (addr_hit[6] & (|(OTP_CTRL_PRIM_PERMIT[6] & ~reg_be))) |
               (addr_hit[7] & (|(OTP_CTRL_PRIM_PERMIT[7] & ~reg_be)))));
  end

  // Generate write-enables
  assign csr0_we = addr_hit[0] & reg_we & !reg_error;

  assign csr0_field0_wd = reg_wdata[0];

  assign csr0_field1_wd = reg_wdata[1];

  assign csr0_field2_wd = reg_wdata[2];

  assign csr0_field3_wd = reg_wdata[13:4];

  assign csr0_field4_wd = reg_wdata[26:16];
  assign csr1_we = addr_hit[1] & reg_we & !reg_error;

  assign csr1_field0_wd = reg_wdata[6:0];

  assign csr1_field1_wd = reg_wdata[7];

  assign csr1_field2_wd = reg_wdata[14:8];

  assign csr1_field3_wd = reg_wdata[15];

  assign csr1_field4_wd = reg_wdata[31:16];
  assign csr2_we = addr_hit[2] & reg_we & !reg_error;

  assign csr2_wd = reg_wdata[0];
  assign csr3_we = addr_hit[3] & reg_we & !reg_error;

  assign csr3_field0_wd = reg_wdata[2:0];

  assign csr3_field1_wd = reg_wdata[13:4];

  assign csr3_field2_wd = reg_wdata[16];
  assign csr4_we = addr_hit[4] & reg_we & !reg_error;

  assign csr4_field0_wd = reg_wdata[9:0];

  assign csr4_field1_wd = reg_wdata[12];

  assign csr4_field2_wd = reg_wdata[13];

  assign csr4_field3_wd = reg_wdata[14];
  assign csr5_we = addr_hit[5] & reg_we & !reg_error;

  assign csr5_field0_wd = reg_wdata[5:0];

  assign csr5_field1_wd = reg_wdata[7:6];

  assign csr5_field6_wd = reg_wdata[31:16];
  assign csr6_we = addr_hit[6] & reg_we & !reg_error;

  assign csr6_field0_wd = reg_wdata[9:0];

  assign csr6_field1_wd = reg_wdata[11];

  assign csr6_field2_wd = reg_wdata[12];

  assign csr6_field3_wd = reg_wdata[31:16];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = csr0_we;
    reg_we_check[1] = csr1_we;
    reg_we_check[2] = csr2_we;
    reg_we_check[3] = csr3_we;
    reg_we_check[4] = csr4_we;
    reg_we_check[5] = csr5_we;
    reg_we_check[6] = csr6_we;
    reg_we_check[7] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = csr0_field0_qs;
        reg_rdata_next[1] = csr0_field1_qs;
        reg_rdata_next[2] = csr0_field2_qs;
        reg_rdata_next[13:4] = csr0_field3_qs;
        reg_rdata_next[26:16] = csr0_field4_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[6:0] = csr1_field0_qs;
        reg_rdata_next[7] = csr1_field1_qs;
        reg_rdata_next[14:8] = csr1_field2_qs;
        reg_rdata_next[15] = csr1_field3_qs;
        reg_rdata_next[31:16] = csr1_field4_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = csr2_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[2:0] = csr3_field0_qs;
        reg_rdata_next[13:4] = csr3_field1_qs;
        reg_rdata_next[16] = csr3_field2_qs;
        reg_rdata_next[17] = csr3_field3_qs;
        reg_rdata_next[18] = csr3_field4_qs;
        reg_rdata_next[19] = csr3_field5_qs;
        reg_rdata_next[20] = csr3_field6_qs;
        reg_rdata_next[21] = csr3_field7_qs;
        reg_rdata_next[22] = csr3_field8_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[9:0] = csr4_field0_qs;
        reg_rdata_next[12] = csr4_field1_qs;
        reg_rdata_next[13] = csr4_field2_qs;
        reg_rdata_next[14] = csr4_field3_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[5:0] = csr5_field0_qs;
        reg_rdata_next[7:6] = csr5_field1_qs;
        reg_rdata_next[8] = csr5_field2_qs;
        reg_rdata_next[11:9] = csr5_field3_qs;
        reg_rdata_next[12] = csr5_field4_qs;
        reg_rdata_next[13] = csr5_field5_qs;
        reg_rdata_next[31:16] = csr5_field6_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[9:0] = csr6_field0_qs;
        reg_rdata_next[11] = csr6_field1_qs;
        reg_rdata_next[12] = csr6_field2_qs;
        reg_rdata_next[31:16] = csr6_field3_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[5:0] = csr7_field0_qs;
        reg_rdata_next[10:8] = csr7_field1_qs;
        reg_rdata_next[14] = csr7_field2_qs;
        reg_rdata_next[15] = csr7_field3_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `CALIPTRA_ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `CALIPTRA_ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `CALIPTRA_ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `CALIPTRA_ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule
