// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef FC_ACCESS_CONTROL_TABLE_SV
`define FC_ACCESS_CONTROL_TABLE_SV

`include "caliptra_ss_includes.svh"
//------------------------------------------------------------------------------
// Generated access control table
// DO NOT EDIT: This file is generated by fc_access_control_table.py
//------------------------------------------------------------------------------

typedef struct packed {
  logic [31:0] lower_addr;  // Lower bound of the address range
  logic [31:0] upper_addr;  // Upper bound of the address range
  logic [3:0]  axi_user_id; // AXI user ID allowed to write
} access_control_entry_t;

localparam int FC_TABLE_NUM_RANGES = 2;

localparam access_control_entry_t access_control_table [FC_TABLE_NUM_RANGES] = '{
  '{ lower_addr: 32'h00000000, upper_addr: 32'h00000080, axi_user_id: CPTRA_SS_STRAP_CLPTRA_CORE_AXI_USER },
  '{ lower_addr: 32'h00000088, upper_addr: 32'h000007A0, axi_user_id: CPTRA_SS_STRAP_MCU_LSU_AXI_USER }
};

`endif // FC_ACCESS_CONTROL_TABLE_SV
