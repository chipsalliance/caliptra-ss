`ifndef aaxi_pkg_caliptra_test_sv
`define aaxi_pkg_caliptra_test_sv

package aaxi_pkg_caliptra_test;

    //`include "aaxi_pkg.sv"
    //`include "aaxi_pkg_test.sv"
    //``include "aaxi_test_caliptra_ss.svh"

endpackage

`endif

